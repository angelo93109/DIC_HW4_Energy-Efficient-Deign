.SUBCKT Convolution_example VSS VDD clk rst_n in_valid In_IFM_1[3] In_IFM_1[2] In_IFM_1[1] In_IFM_1[0] In_IFM_2[3] In_IFM_2[2] In_IFM_2[1] In_IFM_2[0] In_IFM_3[3] In_IFM_3[2] In_IFM_3[1] In_IFM_3[0] In_IFM_4[3] In_IFM_4[2] In_IFM_4[1] In_IFM_4[0] In_Weight_1[3] In_Weight_1[2] In_Weight_1[1] In_Weight_1[0] In_Weight_2[3] In_Weight_2[2] In_Weight_2[1] In_Weight_2[0] In_Weight_3[3] In_Weight_3[2] In_Weight_3[1] In_Weight_3[0] In_Weight_4[3] In_Weight_4[2] In_Weight_4[1] In_Weight_4[0] out_valid Out_OFM[11] Out_OFM[10] Out_OFM[9] Out_OFM[8] Out_OFM[7] Out_OFM[6] Out_OFM[5] Out_OFM[4] Out_OFM[3] Out_OFM[2] Out_OFM[1] Out_OFM[0] 
Xcstate_reg_0_ VSS VDD  n150 clk n162 n253 n116 ASYNC_DFFHx1_ASAP7_75t_R
Xcstate_reg_1_ VSS VDD  n149 clk n162 n182 n115 ASYNC_DFFHx1_ASAP7_75t_R
XIn_4_reg_3_ VSS VDD  n148 clk n162 n178 n114 ASYNC_DFFHx1_ASAP7_75t_R
XIn_4_reg_2_ VSS VDD  n147 clk n162 n176 n113 ASYNC_DFFHx1_ASAP7_75t_R
XIn_4_reg_1_ VSS VDD  n146 clk n162 n151 n112 ASYNC_DFFHx1_ASAP7_75t_R
XIn_4_reg_0_ VSS VDD  n145 clk n162 n171 n111 ASYNC_DFFHx1_ASAP7_75t_R
XIn_1_reg_3_ VSS VDD  n144 clk n162 n208 n110 ASYNC_DFFHx1_ASAP7_75t_R
XIn_1_reg_2_ VSS VDD  n143 clk n162 n254 n109 ASYNC_DFFHx1_ASAP7_75t_R
XIn_1_reg_1_ VSS VDD  n142 clk n162 n200 n108 ASYNC_DFFHx1_ASAP7_75t_R
XIn_1_reg_0_ VSS VDD  n141 clk n162 n188 n107 ASYNC_DFFHx1_ASAP7_75t_R
XIn_2_reg_3_ VSS VDD  n140 clk n162 n186 n106 ASYNC_DFFHx1_ASAP7_75t_R
XIn_2_reg_2_ VSS VDD  n139 clk n162 n179 n105 ASYNC_DFFHx1_ASAP7_75t_R
XIn_2_reg_1_ VSS VDD  n138 clk n162 n210 n104 ASYNC_DFFHx1_ASAP7_75t_R
XIn_2_reg_0_ VSS VDD  n137 clk n162 n194 n103 ASYNC_DFFHx1_ASAP7_75t_R
XIn_3_reg_3_ VSS VDD  n136 clk n162 n193 n102 ASYNC_DFFHx1_ASAP7_75t_R
XIn_3_reg_2_ VSS VDD  n135 clk n162 n195 n101 ASYNC_DFFHx1_ASAP7_75t_R
XIn_3_reg_1_ VSS VDD  n134 clk n162 n198 n100 ASYNC_DFFHx1_ASAP7_75t_R
XIn_3_reg_0_ VSS VDD  n133 clk n162 n229 n99 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts4_reg_3_ VSS VDD  n132 clk n162 n203 n98 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts4_reg_2_ VSS VDD  n131 clk n162 n180 n97 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts4_reg_1_ VSS VDD  n130 clk n162 n233 n96 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts4_reg_0_ VSS VDD  n129 clk n162 n168 n95 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts1_reg_3_ VSS VDD  n128 clk n162 n221 n94 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts1_reg_2_ VSS VDD  n127 clk n162 n201 n93 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts1_reg_1_ VSS VDD  n126 clk n162 n183 n92 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts1_reg_0_ VSS VDD  n125 clk n162 n177 n91 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts2_reg_3_ VSS VDD  n124 clk n162 n191 n90 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts2_reg_2_ VSS VDD  n123 clk n162 n206 n89 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts2_reg_1_ VSS VDD  n122 clk n162 n192 n88 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts2_reg_0_ VSS VDD  n121 clk n162 n174 n87 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts3_reg_3_ VSS VDD  n120 clk n162 n202 n86 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts3_reg_2_ VSS VDD  n119 clk n162 n184 n85 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts3_reg_1_ VSS VDD  n118 clk n162 n196 n84 ASYNC_DFFHx1_ASAP7_75t_R
Xweigts3_reg_0_ VSS VDD  n117 clk n162 n173 n83 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_9_ VSS VDD  n114 clk n162 n209 n81 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_8_ VSS VDD  n113 clk n162 n185 n80 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_7_ VSS VDD  n112 clk n162 n172 n79 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_6_ VSS VDD  n111 clk n162 n197 n78 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_5_ VSS VDD  n110 clk n162 n228 n77 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_4_ VSS VDD  n109 clk n162 n181 n76 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_3_ VSS VDD  n108 clk n162 n175 n75 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_2_ VSS VDD  n107 clk n162 n207 n74 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_1_ VSS VDD  n106 clk n162 n169 n73 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_0_ VSS VDD  n105 clk n162 n187 n72 ASYNC_DFFHx1_ASAP7_75t_R
Xout_valid_reg VSS VDD  n166 clk n162 n170 n70 ASYNC_DFFHx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U128 VSS VDD  DP_OP_20J1_122_6644_n203 DP_OP_20J1_122_6644_n206 DP_OP_20J1_122_6644_n227 DP_OP_20J1_122_6644_n162 DP_OP_20J1_122_6644_n163 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U127 VSS VDD  DP_OP_20J1_122_6644_n230 DP_OP_20J1_122_6644_n254 DP_OP_20J1_122_6644_n251 DP_OP_20J1_122_6644_n160 DP_OP_20J1_122_6644_n161 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U125 VSS VDD  DP_OP_20J1_122_6644_n165 DP_OP_20J1_122_6644_n166 DP_OP_20J1_122_6644_n157 DP_OP_20J1_122_6644_n158 DP_OP_20J1_122_6644_n159 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U122 VSS VDD  DP_OP_20J1_122_6644_n175 DP_OP_20J1_122_6644_n178 DP_OP_20J1_122_6644_n181 DP_OP_20J1_122_6644_n153 DP_OP_20J1_122_6644_n154 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U121 VSS VDD  DP_OP_20J1_122_6644_n199 DP_OP_20J1_122_6644_n202 DP_OP_20J1_122_6644_n205 DP_OP_20J1_122_6644_n151 DP_OP_20J1_122_6644_n152 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U120 VSS VDD  DP_OP_20J1_122_6644_n223 DP_OP_20J1_122_6644_n253 DP_OP_20J1_122_6644_n226 DP_OP_20J1_122_6644_n149 DP_OP_20J1_122_6644_n150 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U119 VSS VDD  DP_OP_20J1_122_6644_n229 DP_OP_20J1_122_6644_n250 DP_OP_20J1_122_6644_n247 DP_OP_20J1_122_6644_n147 DP_OP_20J1_122_6644_n148 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U117 VSS VDD  DP_OP_20J1_122_6644_n162 DP_OP_20J1_122_6644_n144 DP_OP_20J1_122_6644_n160 DP_OP_20J1_122_6644_n145 DP_OP_20J1_122_6644_n146 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U116 VSS VDD  DP_OP_20J1_122_6644_n152 DP_OP_20J1_122_6644_n148 DP_OP_20J1_122_6644_n154 DP_OP_20J1_122_6644_n142 DP_OP_20J1_122_6644_n143 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U114 VSS VDD  DP_OP_20J1_122_6644_n158 DP_OP_20J1_122_6644_n150 DP_OP_20J1_122_6644_n139 DP_OP_20J1_122_6644_n140 DP_OP_20J1_122_6644_n141 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U111 VSS VDD  DP_OP_20J1_122_6644_n177 DP_OP_20J1_122_6644_n180 DP_OP_20J1_122_6644_n195 DP_OP_20J1_122_6644_n135 DP_OP_20J1_122_6644_n136 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U110 VSS VDD  DP_OP_20J1_122_6644_n198 DP_OP_20J1_122_6644_n201 DP_OP_20J1_122_6644_n204 DP_OP_20J1_122_6644_n133 DP_OP_20J1_122_6644_n134 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U109 VSS VDD  DP_OP_20J1_122_6644_n219 DP_OP_20J1_122_6644_n252 DP_OP_20J1_122_6644_n222 DP_OP_20J1_122_6644_n131 DP_OP_20J1_122_6644_n132 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U108 VSS VDD  DP_OP_20J1_122_6644_n225 DP_OP_20J1_122_6644_n249 DP_OP_20J1_122_6644_n228 DP_OP_20J1_122_6644_n129 DP_OP_20J1_122_6644_n130 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U106 VSS VDD  DP_OP_20J1_122_6644_n243 DP_OP_20J1_122_6644_n246 DP_OP_20J1_122_6644_n126 DP_OP_20J1_122_6644_n127 DP_OP_20J1_122_6644_n128 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U104 VSS VDD  DP_OP_20J1_122_6644_n147 DP_OP_20J1_122_6644_n151 DP_OP_20J1_122_6644_n123 DP_OP_20J1_122_6644_n124 DP_OP_20J1_122_6644_n125 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U103 VSS VDD  DP_OP_20J1_122_6644_n132 DP_OP_20J1_122_6644_n149 DP_OP_20J1_122_6644_n130 DP_OP_20J1_122_6644_n121 DP_OP_20J1_122_6644_n122 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U101 VSS VDD  DP_OP_20J1_122_6644_n136 DP_OP_20J1_122_6644_n134 DP_OP_20J1_122_6644_n118 DP_OP_20J1_122_6644_n119 DP_OP_20J1_122_6644_n120 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U99 VSS VDD  DP_OP_20J1_122_6644_n142 DP_OP_20J1_122_6644_n125 DP_OP_20J1_122_6644_n115 DP_OP_20J1_122_6644_n116 DP_OP_20J1_122_6644_n117 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U98 VSS VDD  DP_OP_20J1_122_6644_n120 DP_OP_20J1_122_6644_n122 DP_OP_20J1_122_6644_n140 DP_OP_20J1_122_6644_n113 DP_OP_20J1_122_6644_n114 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U93 VSS VDD  DP_OP_20J1_122_6644_n176 DP_OP_20J1_122_6644_n248 DP_OP_20J1_122_6644_n194 DP_OP_20J1_122_6644_n107 DP_OP_20J1_122_6644_n108 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U92 VSS VDD  DP_OP_20J1_122_6644_n197 DP_OP_20J1_122_6644_n245 DP_OP_20J1_122_6644_n200 DP_OP_20J1_122_6644_n105 DP_OP_20J1_122_6644_n106 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U91 VSS VDD  DP_OP_20J1_122_6644_n218 DP_OP_20J1_122_6644_n242 DP_OP_20J1_122_6644_n221 DP_OP_20J1_122_6644_n103 DP_OP_20J1_122_6644_n104 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U89 VSS VDD  DP_OP_20J1_122_6644_n137 DP_OP_20J1_122_6644_n224 DP_OP_20J1_122_6644_n100 DP_OP_20J1_122_6644_n101 DP_OP_20J1_122_6644_n102 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U87 VSS VDD  DP_OP_20J1_122_6644_n129 DP_OP_20J1_122_6644_n133 DP_OP_20J1_122_6644_n97 DP_OP_20J1_122_6644_n98 DP_OP_20J1_122_6644_n99 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U86 VSS VDD  DP_OP_20J1_122_6644_n104 DP_OP_20J1_122_6644_n131 DP_OP_20J1_122_6644_n106 DP_OP_20J1_122_6644_n95 DP_OP_20J1_122_6644_n96 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U84 VSS VDD  DP_OP_20J1_122_6644_n127 DP_OP_20J1_122_6644_n108 DP_OP_20J1_122_6644_n92 DP_OP_20J1_122_6644_n93 DP_OP_20J1_122_6644_n94 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U82 VSS VDD  DP_OP_20J1_122_6644_n99 DP_OP_20J1_122_6644_n121 DP_OP_20J1_122_6644_n89 DP_OP_20J1_122_6644_n90 DP_OP_20J1_122_6644_n91 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U80 VSS VDD  DP_OP_20J1_122_6644_n96 DP_OP_20J1_122_6644_n119 DP_OP_20J1_122_6644_n86 DP_OP_20J1_122_6644_n87 DP_OP_20J1_122_6644_n88 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U78 VSS VDD  DP_OP_20J1_122_6644_n91 DP_OP_20J1_122_6644_n113 DP_OP_20J1_122_6644_n83 DP_OP_20J1_122_6644_n84 DP_OP_20J1_122_6644_n85 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U74 VSS VDD  DP_OP_20J1_122_6644_n172 DP_OP_20J1_122_6644_n241 DP_OP_20J1_122_6644_n193 DP_OP_20J1_122_6644_n78 DP_OP_20J1_122_6644_n79 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U73 VSS VDD  DP_OP_20J1_122_6644_n196 DP_OP_20J1_122_6644_n220 DP_OP_20J1_122_6644_n217 DP_OP_20J1_122_6644_n76 DP_OP_20J1_122_6644_n77 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U71 VSS VDD  DP_OP_20J1_122_6644_n107 DP_OP_20J1_122_6644_n73 DP_OP_20J1_122_6644_n105 DP_OP_20J1_122_6644_n74 DP_OP_20J1_122_6644_n75 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U69 VSS VDD  DP_OP_20J1_122_6644_n70 DP_OP_20J1_122_6644_n103 DP_OP_20J1_122_6644_n77 DP_OP_20J1_122_6644_n71 DP_OP_20J1_122_6644_n72 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U67 VSS VDD  DP_OP_20J1_122_6644_n101 DP_OP_20J1_122_6644_n79 DP_OP_20J1_122_6644_n67 DP_OP_20J1_122_6644_n68 DP_OP_20J1_122_6644_n69 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U66 VSS VDD  DP_OP_20J1_122_6644_n75 DP_OP_20J1_122_6644_n95 DP_OP_20J1_122_6644_n93 DP_OP_20J1_122_6644_n65 DP_OP_20J1_122_6644_n66 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U64 VSS VDD  DP_OP_20J1_122_6644_n69 DP_OP_20J1_122_6644_n72 DP_OP_20J1_122_6644_n62 DP_OP_20J1_122_6644_n63 DP_OP_20J1_122_6644_n64 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U62 VSS VDD  DP_OP_20J1_122_6644_n87 DP_OP_20J1_122_6644_n66 DP_OP_20J1_122_6644_n59 DP_OP_20J1_122_6644_n60 DP_OP_20J1_122_6644_n61 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U58 VSS VDD  DP_OP_20J1_122_6644_n192 DP_OP_20J1_122_6644_n216 DP_OP_20J1_122_6644_n80 DP_OP_20J1_122_6644_n54 DP_OP_20J1_122_6644_n55 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U56 VSS VDD  DP_OP_20J1_122_6644_n76 DP_OP_20J1_122_6644_n78 DP_OP_20J1_122_6644_n51 DP_OP_20J1_122_6644_n52 DP_OP_20J1_122_6644_n53 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U54 VSS VDD  DP_OP_20J1_122_6644_n71 DP_OP_20J1_122_6644_n74 DP_OP_20J1_122_6644_n48 DP_OP_20J1_122_6644_n49 DP_OP_20J1_122_6644_n50 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U52 VSS VDD  DP_OP_20J1_122_6644_n68 DP_OP_20J1_122_6644_n53 DP_OP_20J1_122_6644_n45 DP_OP_20J1_122_6644_n46 DP_OP_20J1_122_6644_n47 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U51 VSS VDD  DP_OP_20J1_122_6644_n63 DP_OP_20J1_122_6644_n50 DP_OP_20J1_122_6644_n47 DP_OP_20J1_122_6644_n43 DP_OP_20J1_122_6644_n44 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U49 VSS VDD  DP_OP_20J1_122_6644_n52 DP_OP_20J1_122_6644_n56 DP_OP_20J1_122_6644_n40 DP_OP_20J1_122_6644_n41 DP_OP_20J1_122_6644_n42 FAx1_ASAP7_75t_R
XDP_OP_20J1_122_6644_U48 VSS VDD  DP_OP_20J1_122_6644_n42 DP_OP_20J1_122_6644_n49 DP_OP_20J1_122_6644_n46 DP_OP_20J1_122_6644_n38 DP_OP_20J1_122_6644_n39 FAx1_ASAP7_75t_R
XU163 VSS VDD  n369 n160 n370 XNOR2xp5_ASAP7_75t_R
XU164 VSS VDD  DP_OP_20J1_122_6644_n143 n363 n361 XOR2xp5_ASAP7_75t_R
XU165 VSS VDD  n160 n238 INVx2_ASAP7_75t_R
XU166 VSS VDD  n159 n239 INVx2_ASAP7_75t_R
XU167 VSS VDD  n227 n345 INVx3_ASAP7_75t_R
XU168 VSS VDD  n152 n343 INVx2_ASAP7_75t_R
XU169 VSS VDD  n241 n344 INVx2_ASAP7_75t_R
XU170 VSS VDD  n252 n297 INVx3_ASAP7_75t_R
XU171 VSS VDD  n226 n251 INVx3_ASAP7_75t_R
XU172 VSS VDD  n222 n281 INVx2_ASAP7_75t_R
XU173 VSS VDD  n101 n157 BUFx5_ASAP7_75t_R
XU174 VSS VDD  n103 n156 BUFx5_ASAP7_75t_R
XU175 VSS VDD  n83 n158 BUFx5_ASAP7_75t_R
XU176 VSS VDD  n98 n154 BUFx5_ASAP7_75t_R
XU177 VSS VDD  n86 n155 BUFx5_ASAP7_75t_R
XU178 VSS VDD  n87 n161 BUFx5_ASAP7_75t_R
XU179 VSS VDD  n102 n153 BUFx5_ASAP7_75t_R
XU180 VSS VDD  n111 n152 BUFx5_ASAP7_75t_R
XU181 VSS VDD  n110 n214 BUFx5_ASAP7_75t_R
XU182 VSS VDD  n115 n383 BUFx5_ASAP7_75t_R
XU183 VSS VDD  n116 n385 BUFx5_ASAP7_75t_R
XU184 VSS VDD  n109 n213 BUFx5_ASAP7_75t_R
XU185 VSS VDD  n108 n212 BUFx5_ASAP7_75t_R
XU186 VSS VDD  n107 n220 BUFx5_ASAP7_75t_R
XU187 VSS VDD  n106 n218 BUFx5_ASAP7_75t_R
XU188 VSS VDD  n104 n216 BUFx5_ASAP7_75t_R
XU189 VSS VDD  n94 n243 BUFx5_ASAP7_75t_R
XU190 VSS VDD  n105 n217 BUFx5_ASAP7_75t_R
XU191 VSS VDD  n100 n225 BUFx5_ASAP7_75t_R
XU192 VSS VDD  n90 n246 BUFx5_ASAP7_75t_R
XU193 VSS VDD  n91 n242 BUFx5_ASAP7_75t_R
XU194 VSS VDD  n92 n245 BUFx5_ASAP7_75t_R
XU195 VSS VDD  n93 n244 BUFx5_ASAP7_75t_R
XU196 VSS VDD  n89 n247 BUFx5_ASAP7_75t_R
XU197 VSS VDD  n88 n248 BUFx5_ASAP7_75t_R
XU198 VSS VDD  n84 n250 BUFx5_ASAP7_75t_R
XU199 VSS VDD  n85 n249 BUFx5_ASAP7_75t_R
XU200 VSS VDD  n114 n252 BUFx8_ASAP7_75t_R
XU201 VSS VDD  n167 n370 N110 NOR2xp33_ASAP7_75t_R
XU202 VSS VDD  n286 n285 n147 NAND2xp33_ASAP7_75t_R
XU203 VSS VDD  n268 n267 n136 NAND2xp33_ASAP7_75t_R
XU204 VSS VDD  n259 n258 n137 NAND2xp33_ASAP7_75t_R
XU205 VSS VDD  n294 n293 n146 NAND2xp33_ASAP7_75t_R
XU206 VSS VDD  n283 n282 n131 NAND2xp33_ASAP7_75t_R
XU207 VSS VDD  n273 n272 n133 NAND2xp33_ASAP7_75t_R
XU208 VSS VDD  n277 n276 n135 NAND2xp33_ASAP7_75t_R
XU209 VSS VDD  n305 n304 n121 NAND2xp33_ASAP7_75t_R
XU210 VSS VDD  n264 n263 n130 NAND2xp33_ASAP7_75t_R
XU211 VSS VDD  n340 n339 n117 NAND2xp33_ASAP7_75t_R
XU212 VSS VDD  n314 n313 n140 NAND2xp33_ASAP7_75t_R
XU213 VSS VDD  n321 n320 n141 NAND2xp33_ASAP7_75t_R
XU214 VSS VDD  n329 n328 n142 NAND2xp33_ASAP7_75t_R
XU215 VSS VDD  n338 n337 n143 NAND2xp33_ASAP7_75t_R
XU216 VSS VDD  n292 n291 n128 NAND2xp33_ASAP7_75t_R
XU217 VSS VDD  n262 n261 n134 NAND2xp33_ASAP7_75t_R
XU218 VSS VDD  n296 n295 n138 NAND2xp33_ASAP7_75t_R
XU219 VSS VDD  n311 n310 n139 NAND2xp33_ASAP7_75t_R
XU220 VSS VDD  n302 n301 n124 NAND2xp33_ASAP7_75t_R
XU221 VSS VDD  n332 n331 n125 NAND2xp33_ASAP7_75t_R
XU222 VSS VDD  n280 n279 n126 NAND2xp33_ASAP7_75t_R
XU223 VSS VDD  n271 n270 n127 NAND2xp33_ASAP7_75t_R
XU224 VSS VDD  n299 n298 n148 NAND2xp33_ASAP7_75t_R
XU225 VSS VDD  n324 n323 n119 NAND2xp33_ASAP7_75t_R
XU226 VSS VDD  n327 n326 n122 NAND2xp33_ASAP7_75t_R
XU227 VSS VDD  n317 n316 n123 NAND2xp33_ASAP7_75t_R
XU228 VSS VDD  n335 n334 n118 NAND2xp33_ASAP7_75t_R
XU229 VSS VDD  n308 n307 n120 NAND2xp33_ASAP7_75t_R
XU230 VSS VDD  n266 n265 n132 NAND2xp33_ASAP7_75t_R
XU231 VSS VDD  n112 n241 BUFx5_ASAP7_75t_R
XU232 VSS VDD  n275 n274 n145 NAND2xp33_ASAP7_75t_R
XU233 VSS VDD  n95 n227 BUFx5_ASAP7_75t_R
XU234 VSS VDD  n97 n222 BUFx5_ASAP7_75t_R
XU235 VSS VDD  n223 n284 INVx3_ASAP7_75t_R
XU236 VSS VDD  n113 n223 BUFx5_ASAP7_75t_R
XU237 VSS VDD  n99 n236 BUFx5_ASAP7_75t_R
XU238 VSS VDD  DP_OP_20J1_122_6644_n88 n159 BUFx4_ASAP7_75t_R
XU239 VSS VDD  DP_OP_20J1_122_6644_n61 n160 BUFx4_ASAP7_75t_R
XU240 VSS VDD  n256 n255 n257 NAND2xp33_ASAP7_75t_R
XU241 VSS VDD  DP_OP_20J1_122_6644_n73 n257 DP_OP_20J1_122_6644_n97 NAND2xp33_ASAP7_75t_R
XU242 VSS VDD  DP_OP_20J1_122_6644_n166 n354 n357 NOR2xp33_ASAP7_75t_R
XU243 VSS VDD  In_Weight_2[0] in_valid n305 NAND2xp33_ASAP7_75t_R
XU244 VSS VDD  in_valid In_Weight_1[3] n292 NAND2xp33_ASAP7_75t_R
XU245 VSS VDD  in_valid In_IFM_3[3] n268 NAND2xp33_ASAP7_75t_R
XU246 VSS VDD  in_valid In_IFM_1[2] n338 NAND2xp33_ASAP7_75t_R
XU247 VSS VDD  n319 n318 n129 NAND2xp33_ASAP7_75t_R
XU248 VSS VDD  n289 n288 n144 NAND2xp33_ASAP7_75t_R
XU249 VSS VDD  in_valid n386 n260 NOR2x1_ASAP7_75t_R
XU250 VSS VDD  In_Weight_3[0] in_valid n340 NAND2xp5_ASAP7_75t_R
XU251 VSS VDD  in_valid In_IFM_4[1] n294 NAND2xp5_ASAP7_75t_R
XU252 VSS VDD  in_valid In_IFM_3[1] n262 NAND2xp5_ASAP7_75t_R
XU253 VSS VDD  in_valid In_Weight_3[2] n324 NAND2xp5_ASAP7_75t_R
XU254 VSS VDD  in_valid In_Weight_3[3] n308 NAND2xp5_ASAP7_75t_R
XU255 VSS VDD  In_IFM_4[0] in_valid n275 NAND2xp5_ASAP7_75t_R
XU256 VSS VDD  in_valid In_Weight_4[3] n266 NAND2xp5_ASAP7_75t_R
XU257 VSS VDD  in_valid In_Weight_1[2] n271 NAND2xp5_ASAP7_75t_R
XU258 VSS VDD  in_valid In_IFM_4[2] n286 NAND2xp5_ASAP7_75t_R
XU259 VSS VDD  in_valid In_IFM_3[2] n277 NAND2xp5_ASAP7_75t_R
XU260 VSS VDD  in_valid In_IFM_4[3] n299 NAND2xp5_ASAP7_75t_R
XU261 VSS VDD  in_valid In_IFM_1[3] n289 NAND2xp5_ASAP7_75t_R
XU262 VSS VDD  in_valid In_Weight_3[1] n335 NAND2xp5_ASAP7_75t_R
XU263 VSS VDD  in_valid In_IFM_1[1] n329 NAND2xp5_ASAP7_75t_R
XU264 VSS VDD  In_IFM_3[0] in_valid n273 NAND2xp5_ASAP7_75t_R
XU265 VSS VDD  In_Weight_1[0] in_valid n332 NAND2xp5_ASAP7_75t_R
XU266 VSS VDD  in_valid In_Weight_4[1] n264 NAND2xp5_ASAP7_75t_R
XU267 VSS VDD  In_IFM_2[0] in_valid n259 NAND2xp5_ASAP7_75t_R
XU268 VSS VDD  in_valid In_IFM_2[1] n296 NAND2xp5_ASAP7_75t_R
XU269 VSS VDD  in_valid In_Weight_2[3] n302 NAND2xp5_ASAP7_75t_R
XU270 VSS VDD  in_valid In_IFM_2[2] n311 NAND2xp5_ASAP7_75t_R
XU271 VSS VDD  in_valid In_IFM_2[3] n314 NAND2xp5_ASAP7_75t_R
XU272 VSS VDD  in_valid In_Weight_2[2] n317 NAND2xp5_ASAP7_75t_R
XU273 VSS VDD  in_valid In_Weight_4[2] n283 NAND2xp5_ASAP7_75t_R
XU274 VSS VDD  in_valid In_Weight_1[1] n280 NAND2xp5_ASAP7_75t_R
XU275 VSS VDD  in_valid In_Weight_2[1] n327 NAND2xp5_ASAP7_75t_R
XU276 VSS VDD  In_Weight_4[0] in_valid n319 NAND2xp5_ASAP7_75t_R
XU277 VSS VDD  In_IFM_1[0] in_valid n321 NAND2xp5_ASAP7_75t_R
XU278 VSS VDD  DP_OP_20J1_122_6644_n38 n380 INVxp67_ASAP7_75t_R
XU279 VSS VDD  n236 n235 INVx1_ASAP7_75t_R
XU280 VSS VDD  n158 n232 INVx1_ASAP7_75t_R
XU281 VSS VDD  n156 n231 INVx1_ASAP7_75t_R
XU282 VSS VDD  n157 n237 INVx1_ASAP7_75t_R
XU283 VSS VDD  n155 n306 INVx1_ASAP7_75t_R
XU284 VSS VDD  n385 n204 INVx2_ASAP7_75t_R
XU285 VSS VDD  n383 n205 INVx2_ASAP7_75t_R
XU286 VSS VDD  n162 TIELOx1_ASAP7_75t_R
XU287 VSS VDD  n165 TIEHIx1_ASAP7_75t_R
XU288 VSS VDD  n165 Out_OFM[10] INVxp33_ASAP7_75t_R
XU289 VSS VDD  n165 Out_OFM[11] INVxp33_ASAP7_75t_R
XU290 VSS VDD  n161 n303 INVx2_ASAP7_75t_R
XU291 VSS VDD  n154 n234 INVx2_ASAP7_75t_R
XU292 VSS VDD  n153 n230 INVx2_ASAP7_75t_R
XU293 VSS VDD  n220 n219 INVx2_ASAP7_75t_R
XU294 VSS VDD  n216 n215 INVx2_ASAP7_75t_R
XU295 VSS VDD  n212 n211 INVx2_ASAP7_75t_R
XU296 VSS VDD  n225 n224 INVx2_ASAP7_75t_R
XU297 VSS VDD  n383 n385 n166 NOR2xp33_ASAP7_75t_R
XU298 VSS VDD  n383 n385 n167 OR2x2_ASAP7_75t_R
XU299 VSS VDD  rst_n n168 INVx8_ASAP7_75t_R
XU300 VSS VDD  rst_n n169 INVx8_ASAP7_75t_R
XU301 VSS VDD  rst_n n170 INVx8_ASAP7_75t_R
XU302 VSS VDD  rst_n n171 INVx8_ASAP7_75t_R
XU303 VSS VDD  rst_n n172 INVx8_ASAP7_75t_R
XU304 VSS VDD  rst_n n173 INVx8_ASAP7_75t_R
XU305 VSS VDD  rst_n n174 INVx8_ASAP7_75t_R
XU306 VSS VDD  rst_n n175 INVx8_ASAP7_75t_R
XU307 VSS VDD  rst_n n176 INVx8_ASAP7_75t_R
XU308 VSS VDD  rst_n n177 INVx8_ASAP7_75t_R
XU309 VSS VDD  rst_n n178 INVx8_ASAP7_75t_R
XU310 VSS VDD  rst_n n179 INVx8_ASAP7_75t_R
XU311 VSS VDD  rst_n n180 INVx8_ASAP7_75t_R
XU312 VSS VDD  rst_n n181 INVx8_ASAP7_75t_R
XU313 VSS VDD  rst_n n182 INVx8_ASAP7_75t_R
XU314 VSS VDD  rst_n n183 INVx8_ASAP7_75t_R
XU315 VSS VDD  rst_n n184 INVx8_ASAP7_75t_R
XU316 VSS VDD  rst_n n185 INVx8_ASAP7_75t_R
XU317 VSS VDD  rst_n n186 INVx8_ASAP7_75t_R
XU318 VSS VDD  rst_n n187 INVx8_ASAP7_75t_R
XU319 VSS VDD  rst_n n188 INVx8_ASAP7_75t_R
XU320 VSS VDD  n359 n358 n357 n189 MAJIxp5_ASAP7_75t_R
XU321 VSS VDD  DP_OP_20J1_122_6644_n141 DP_OP_20J1_122_6644_n143 n363 n190 MAJIxp5_ASAP7_75t_R
XU322 VSS VDD  rst_n n191 INVx8_ASAP7_75t_R
XU323 VSS VDD  rst_n n192 INVx8_ASAP7_75t_R
XU324 VSS VDD  rst_n n193 INVx8_ASAP7_75t_R
XU325 VSS VDD  rst_n n194 INVx8_ASAP7_75t_R
XU326 VSS VDD  rst_n n195 INVx8_ASAP7_75t_R
XU327 VSS VDD  rst_n n196 INVx8_ASAP7_75t_R
XU328 VSS VDD  rst_n n197 INVx8_ASAP7_75t_R
XU329 VSS VDD  rst_n n198 INVx8_ASAP7_75t_R
XU330 VSS VDD  n359 n358 n357 n199 MAJx2_ASAP7_75t_R
XU331 VSS VDD  rst_n n200 INVx8_ASAP7_75t_R
XU332 VSS VDD  rst_n n201 INVx8_ASAP7_75t_R
XU333 VSS VDD  rst_n n202 INVx8_ASAP7_75t_R
XU334 VSS VDD  rst_n n203 INVx8_ASAP7_75t_R
XU335 VSS VDD  n96 n226 BUFx5_ASAP7_75t_R
XU336 VSS VDD  n217 n309 INVx2_ASAP7_75t_R
XU337 VSS VDD  n218 n312 INVx2_ASAP7_75t_R
XU338 VSS VDD  n213 n336 INVx2_ASAP7_75t_R
XU339 VSS VDD  n214 n287 INVx2_ASAP7_75t_R
XU340 VSS VDD  n248 n325 INVx2_ASAP7_75t_R
XU341 VSS VDD  n249 n322 INVx2_ASAP7_75t_R
XU342 VSS VDD  n250 n333 INVx2_ASAP7_75t_R
XU343 VSS VDD  n242 n330 INVx2_ASAP7_75t_R
XU344 VSS VDD  n244 n269 INVx2_ASAP7_75t_R
XU345 VSS VDD  n245 n278 INVx2_ASAP7_75t_R
XU346 VSS VDD  n246 n300 INVx2_ASAP7_75t_R
XU347 VSS VDD  n247 n315 INVx2_ASAP7_75t_R
XU348 VSS VDD  n243 n290 INVx2_ASAP7_75t_R
XU349 VSS VDD  DP_OP_20J1_122_6644_n141 DP_OP_20J1_122_6644_n143 n363 n365 MAJx2_ASAP7_75t_R
XU350 VSS VDD  DP_OP_20J1_122_6644_n146 DP_OP_20J1_122_6644_n139 INVx1_ASAP7_75t_R
XU351 VSS VDD  DP_OP_20J1_122_6644_n135 DP_OP_20J1_122_6644_n100 INVx1_ASAP7_75t_R
XU352 VSS VDD  DP_OP_20J1_122_6644_n153 DP_OP_20J1_122_6644_n126 INVx1_ASAP7_75t_R
XU353 VSS VDD  rst_n n206 INVx8_ASAP7_75t_R
XU354 VSS VDD  rst_n n207 INVx8_ASAP7_75t_R
XU355 VSS VDD  DP_OP_20J1_122_6644_n90 DP_OP_20J1_122_6644_n62 INVx1_ASAP7_75t_R
XU356 VSS VDD  DP_OP_20J1_122_6644_n65 DP_OP_20J1_122_6644_n45 INVx1_ASAP7_75t_R
XU357 VSS VDD  rst_n n208 INVx8_ASAP7_75t_R
XU358 VSS VDD  DP_OP_20J1_122_6644_n54 DP_OP_20J1_122_6644_n40 INVx1_ASAP7_75t_R
XU359 VSS VDD  DP_OP_20J1_122_6644_n55 DP_OP_20J1_122_6644_n48 INVx1_ASAP7_75t_R
XU360 VSS VDD  rst_n n209 INVx8_ASAP7_75t_R
XU361 VSS VDD  rst_n n210 INVx8_ASAP7_75t_R
XU362 VSS VDD  DP_OP_20J1_122_6644_n116 DP_OP_20J1_122_6644_n86 INVx1_ASAP7_75t_R
XU363 VSS VDD  DP_OP_20J1_122_6644_n84 DP_OP_20J1_122_6644_n59 INVx1_ASAP7_75t_R
XU364 VSS VDD  rst_n n221 INVx8_ASAP7_75t_R
XU365 VSS VDD  rst_n n228 INVx8_ASAP7_75t_R
XU366 VSS VDD  rst_n n229 INVx8_ASAP7_75t_R
XU367 VSS VDD  rst_n n233 INVx8_ASAP7_75t_R
XU368 VSS VDD  DP_OP_20J1_122_6644_n124 DP_OP_20J1_122_6644_n92 INVx1_ASAP7_75t_R
XU369 VSS VDD  DP_OP_20J1_122_6644_n163 DP_OP_20J1_122_6644_n157 INVx1_ASAP7_75t_R
XU370 VSS VDD  DP_OP_20J1_122_6644_n145 DP_OP_20J1_122_6644_n118 INVx1_ASAP7_75t_R
XU371 VSS VDD  DP_OP_20J1_122_6644_n98 DP_OP_20J1_122_6644_n67 INVx1_ASAP7_75t_R
XU372 VSS VDD  DP_OP_20J1_122_6644_n102 DP_OP_20J1_122_6644_n89 INVx1_ASAP7_75t_R
XU373 VSS VDD  DP_OP_20J1_122_6644_n128 DP_OP_20J1_122_6644_n115 INVx1_ASAP7_75t_R
XU374 VSS VDD  DP_OP_20J1_122_6644_n94 DP_OP_20J1_122_6644_n83 INVx1_ASAP7_75t_R
XU375 VSS VDD  DP_OP_20J1_122_6644_n42 DP_OP_20J1_122_6644_n49 DP_OP_20J1_122_6644_n46 n240 MAJIxp5_ASAP7_75t_R
XU376 VSS VDD  n240 n378 n379 XNOR2xp5_ASAP7_75t_R
XU377 VSS VDD  rst_n n253 INVx8_ASAP7_75t_R
XU378 VSS VDD  rst_n n254 INVx8_ASAP7_75t_R
XU379 VSS VDD  rst_n n151 INVx8_ASAP7_75t_R
XU380 VSS VDD  n80 Out_OFM[8] INVxp33_ASAP7_75t_R
XU381 VSS VDD  n74 Out_OFM[2] INVxp33_ASAP7_75t_R
XU382 VSS VDD  n77 Out_OFM[5] INVxp33_ASAP7_75t_R
XU383 VSS VDD  n75 Out_OFM[3] INVxp33_ASAP7_75t_R
XU384 VSS VDD  n81 Out_OFM[9] INVxp33_ASAP7_75t_R
XU385 VSS VDD  n70 out_valid INVxp33_ASAP7_75t_R
XU386 VSS VDD  n72 Out_OFM[0] INVxp33_ASAP7_75t_R
XU387 VSS VDD  n79 Out_OFM[7] INVxp33_ASAP7_75t_R
XU388 VSS VDD  n76 Out_OFM[4] INVxp33_ASAP7_75t_R
XU389 VSS VDD  n78 Out_OFM[6] INVxp33_ASAP7_75t_R
XU390 VSS VDD  n73 Out_OFM[1] INVxp33_ASAP7_75t_R
XU391 VSS VDD  n297 n284 n251 n281 DP_OP_20J1_122_6644_n73 NAND4xp25_ASAP7_75t_R
XU392 VSS VDD  n251 n297 n256 NAND2xp33_ASAP7_75t_R
XU393 VSS VDD  n284 n281 n255 NAND2xp33_ASAP7_75t_R
XU394 VSS VDD  n204 n205 n386 NOR2xp33_ASAP7_75t_R
XU395 VSS VDD  n231 n260 n258 NAND2xp33_ASAP7_75t_R
XU396 VSS VDD  n224 n260 n261 NAND2xp33_ASAP7_75t_R
XU397 VSS VDD  n251 n260 n263 NAND2xp33_ASAP7_75t_R
XU398 VSS VDD  n234 n260 n265 NAND2xp33_ASAP7_75t_R
XU399 VSS VDD  n230 n260 n267 NAND2xp33_ASAP7_75t_R
XU400 VSS VDD  n269 n260 n270 NAND2xp33_ASAP7_75t_R
XU401 VSS VDD  n235 n260 n272 NAND2xp33_ASAP7_75t_R
XU402 VSS VDD  n343 n260 n274 NAND2xp33_ASAP7_75t_R
XU403 VSS VDD  n237 n260 n276 NAND2xp33_ASAP7_75t_R
XU404 VSS VDD  n278 n260 n279 NAND2xp33_ASAP7_75t_R
XU405 VSS VDD  n281 n260 n282 NAND2xp33_ASAP7_75t_R
XU406 VSS VDD  n284 n260 n285 NAND2xp33_ASAP7_75t_R
XU407 VSS VDD  n287 n260 n288 NAND2xp33_ASAP7_75t_R
XU408 VSS VDD  n290 n260 n291 NAND2xp33_ASAP7_75t_R
XU409 VSS VDD  n344 n260 n293 NAND2xp33_ASAP7_75t_R
XU410 VSS VDD  n215 n260 n295 NAND2xp33_ASAP7_75t_R
XU411 VSS VDD  n297 n260 n298 NAND2xp33_ASAP7_75t_R
XU412 VSS VDD  n300 n260 n301 NAND2xp33_ASAP7_75t_R
XU413 VSS VDD  n260 n303 n304 NAND2xp33_ASAP7_75t_R
XU414 VSS VDD  n306 n260 n307 NAND2xp33_ASAP7_75t_R
XU415 VSS VDD  n309 n260 n310 NAND2xp33_ASAP7_75t_R
XU416 VSS VDD  n312 n260 n313 NAND2xp33_ASAP7_75t_R
XU417 VSS VDD  n315 n260 n316 NAND2xp33_ASAP7_75t_R
XU418 VSS VDD  n345 n260 n318 NAND2xp33_ASAP7_75t_R
XU419 VSS VDD  n219 n260 n320 NAND2xp33_ASAP7_75t_R
XU420 VSS VDD  n322 n260 n323 NAND2xp33_ASAP7_75t_R
XU421 VSS VDD  n325 n260 n326 NAND2xp33_ASAP7_75t_R
XU422 VSS VDD  n211 n260 n328 NAND2xp33_ASAP7_75t_R
XU423 VSS VDD  n330 n260 n331 NAND2xp33_ASAP7_75t_R
XU424 VSS VDD  n333 n260 n334 NAND2xp33_ASAP7_75t_R
XU425 VSS VDD  n336 n260 n337 NAND2xp33_ASAP7_75t_R
XU426 VSS VDD  n232 n260 n339 NAND2xp33_ASAP7_75t_R
XU427 VSS VDD  n227 n252 n342 NOR2xp33_ASAP7_75t_R
XU428 VSS VDD  n223 n226 n341 NOR2xp33_ASAP7_75t_R
XU429 VSS VDD  n342 n341 A0  DP_OP_20J1_122_6644_n123 HAxp5_ASAP7_75t_R
XU430 VSS VDD  n252 n227 n223 n226 DP_OP_20J1_122_6644_n137 NOR4xp25_ASAP7_75t_R
XU431 VSS VDD  n345 n343 n344 n251 DP_OP_20J1_122_6644_n144 NAND4xp25_ASAP7_75t_R
XU432 VSS VDD  n152 n226 n347 NOR2xp33_ASAP7_75t_R
XU433 VSS VDD  n345 n344 n346 NAND2xp33_ASAP7_75t_R
XU434 VSS VDD  n347 n346 A1  DP_OP_20J1_122_6644_n165 HAxp5_ASAP7_75t_R
XU435 VSS VDD  n161 n156 n158 n236 DP_OP_20J1_122_6644_n166 NOR4xp25_ASAP7_75t_R
XU436 VSS VDD  n154 n223 DP_OP_20J1_122_6644_n172 NOR2xp33_ASAP7_75t_R
XU437 VSS VDD  n227 n223 DP_OP_20J1_122_6644_n175 NOR2xp33_ASAP7_75t_R
XU438 VSS VDD  n241 n154 DP_OP_20J1_122_6644_n176 NOR2xp33_ASAP7_75t_R
XU439 VSS VDD  n241 n222 DP_OP_20J1_122_6644_n177 NOR2xp33_ASAP7_75t_R
XU440 VSS VDD  n241 n226 DP_OP_20J1_122_6644_n178 NOR2xp33_ASAP7_75t_R
XU441 VSS VDD  n152 n154 DP_OP_20J1_122_6644_n180 NOR2xp33_ASAP7_75t_R
XU442 VSS VDD  n152 n222 DP_OP_20J1_122_6644_n181 NOR2xp33_ASAP7_75t_R
XU443 VSS VDD  n218 n246 DP_OP_20J1_122_6644_n192 NOR2xp33_ASAP7_75t_R
XU444 VSS VDD  n218 n247 DP_OP_20J1_122_6644_n193 NOR2xp33_ASAP7_75t_R
XU445 VSS VDD  n218 n248 DP_OP_20J1_122_6644_n194 NOR2xp33_ASAP7_75t_R
XU446 VSS VDD  n218 n161 DP_OP_20J1_122_6644_n195 NOR2xp33_ASAP7_75t_R
XU447 VSS VDD  n217 n246 DP_OP_20J1_122_6644_n196 NOR2xp33_ASAP7_75t_R
XU448 VSS VDD  n217 n247 DP_OP_20J1_122_6644_n197 NOR2xp33_ASAP7_75t_R
XU449 VSS VDD  n217 n248 DP_OP_20J1_122_6644_n198 NOR2xp33_ASAP7_75t_R
XU450 VSS VDD  n217 n161 DP_OP_20J1_122_6644_n199 NOR2xp33_ASAP7_75t_R
XU451 VSS VDD  n216 n246 DP_OP_20J1_122_6644_n200 NOR2xp33_ASAP7_75t_R
XU452 VSS VDD  n216 n247 DP_OP_20J1_122_6644_n201 NOR2xp33_ASAP7_75t_R
XU453 VSS VDD  n216 n248 DP_OP_20J1_122_6644_n202 NOR2xp33_ASAP7_75t_R
XU454 VSS VDD  n216 n161 DP_OP_20J1_122_6644_n203 NOR2xp33_ASAP7_75t_R
XU455 VSS VDD  n246 n156 DP_OP_20J1_122_6644_n204 NOR2xp33_ASAP7_75t_R
XU456 VSS VDD  n247 n156 DP_OP_20J1_122_6644_n205 NOR2xp33_ASAP7_75t_R
XU457 VSS VDD  n248 n156 DP_OP_20J1_122_6644_n206 NOR2xp33_ASAP7_75t_R
XU458 VSS VDD  n214 n243 DP_OP_20J1_122_6644_n216 NOR2xp33_ASAP7_75t_R
XU459 VSS VDD  n214 n244 DP_OP_20J1_122_6644_n217 NOR2xp33_ASAP7_75t_R
XU460 VSS VDD  n214 n245 DP_OP_20J1_122_6644_n218 NOR2xp33_ASAP7_75t_R
XU461 VSS VDD  n214 n242 DP_OP_20J1_122_6644_n219 NOR2xp33_ASAP7_75t_R
XU462 VSS VDD  n213 n243 DP_OP_20J1_122_6644_n220 NOR2xp33_ASAP7_75t_R
XU463 VSS VDD  n213 n244 DP_OP_20J1_122_6644_n221 NOR2xp33_ASAP7_75t_R
XU464 VSS VDD  n213 n245 DP_OP_20J1_122_6644_n222 NOR2xp33_ASAP7_75t_R
XU465 VSS VDD  n242 n213 DP_OP_20J1_122_6644_n223 NOR2xp33_ASAP7_75t_R
XU466 VSS VDD  n243 n212 DP_OP_20J1_122_6644_n224 NOR2xp33_ASAP7_75t_R
XU467 VSS VDD  n212 n244 DP_OP_20J1_122_6644_n225 NOR2xp33_ASAP7_75t_R
XU468 VSS VDD  n212 n245 DP_OP_20J1_122_6644_n226 NOR2xp33_ASAP7_75t_R
XU469 VSS VDD  n242 n212 DP_OP_20J1_122_6644_n227 NOR2xp33_ASAP7_75t_R
XU470 VSS VDD  n220 n243 DP_OP_20J1_122_6644_n228 NOR2xp33_ASAP7_75t_R
XU471 VSS VDD  n220 n244 DP_OP_20J1_122_6644_n229 NOR2xp33_ASAP7_75t_R
XU472 VSS VDD  n245 n220 DP_OP_20J1_122_6644_n230 NOR2xp33_ASAP7_75t_R
XU473 VSS VDD  n249 n153 DP_OP_20J1_122_6644_n241 NOR2xp33_ASAP7_75t_R
XU474 VSS VDD  n250 n153 DP_OP_20J1_122_6644_n242 NOR2xp33_ASAP7_75t_R
XU475 VSS VDD  n153 n158 DP_OP_20J1_122_6644_n243 NOR2xp33_ASAP7_75t_R
XU476 VSS VDD  n249 n157 DP_OP_20J1_122_6644_n245 NOR2xp33_ASAP7_75t_R
XU477 VSS VDD  n250 n157 DP_OP_20J1_122_6644_n246 NOR2xp33_ASAP7_75t_R
XU478 VSS VDD  n158 n157 DP_OP_20J1_122_6644_n247 NOR2xp33_ASAP7_75t_R
XU479 VSS VDD  n225 n155 DP_OP_20J1_122_6644_n248 NOR2xp33_ASAP7_75t_R
XU480 VSS VDD  n225 n249 DP_OP_20J1_122_6644_n249 NOR2xp33_ASAP7_75t_R
XU481 VSS VDD  n250 n225 DP_OP_20J1_122_6644_n250 NOR2xp33_ASAP7_75t_R
XU482 VSS VDD  n225 n158 DP_OP_20J1_122_6644_n251 NOR2xp33_ASAP7_75t_R
XU483 VSS VDD  n236 n155 DP_OP_20J1_122_6644_n252 NOR2xp33_ASAP7_75t_R
XU484 VSS VDD  n249 n236 DP_OP_20J1_122_6644_n253 NOR2xp33_ASAP7_75t_R
XU485 VSS VDD  n250 n236 DP_OP_20J1_122_6644_n254 NOR2xp33_ASAP7_75t_R
XU486 VSS VDD  n154 n252 n349 NOR2xp33_ASAP7_75t_R
XU487 VSS VDD  n153 n155 n348 NOR2xp33_ASAP7_75t_R
XU488 VSS VDD  n349 n348 A2  DP_OP_20J1_122_6644_n51 HAxp5_ASAP7_75t_R
XU489 VSS VDD  n252 n153 n154 n155 DP_OP_20J1_122_6644_n56 NOR4xp25_ASAP7_75t_R
XU490 VSS VDD  n252 n222 n351 NOR2xp33_ASAP7_75t_R
XU491 VSS VDD  n157 n155 n350 NOR2xp33_ASAP7_75t_R
XU492 VSS VDD  n351 n350 A3  DP_OP_20J1_122_6644_n70 HAxp5_ASAP7_75t_R
XU493 VSS VDD  n157 n155 n222 n252 DP_OP_20J1_122_6644_n80 NOR4xp25_ASAP7_75t_R
XU494 VSS VDD  n161 n156 n353 NOR2xp33_ASAP7_75t_R
XU495 VSS VDD  n236 n158 n352 NOR2xp33_ASAP7_75t_R
XU496 VSS VDD  n353 n352 n354 NOR2xp33_ASAP7_75t_R
XU497 VSS VDD  n227 n152 n359 NOR2xp33_ASAP7_75t_R
XU498 VSS VDD  n220 n242 n358 NOR2xp33_ASAP7_75t_R
XU499 VSS VDD  n359 n358 n355 XOR2xp5_ASAP7_75t_R
XU500 VSS VDD  n357 n355 A4  n356 HAxp5_ASAP7_75t_R
XU501 VSS VDD  n167 n356 N105 NOR2xp33_ASAP7_75t_R
XU502 VSS VDD  DP_OP_20J1_122_6644_n159 DP_OP_20J1_122_6644_n161 n199 A5  n360 FAx1_ASAP7_75t_R
XU503 VSS VDD  n167 n360 N106 NOR2xp33_ASAP7_75t_R
XU504 VSS VDD  n189 DP_OP_20J1_122_6644_n161 DP_OP_20J1_122_6644_n159 n363 MAJIxp5_ASAP7_75t_R
XU505 VSS VDD  DP_OP_20J1_122_6644_n141 n361 A6  n362 HAxp5_ASAP7_75t_R
XU506 VSS VDD  n167 n362 N107 NOR2xp33_ASAP7_75t_R
XU507 VSS VDD  DP_OP_20J1_122_6644_n114 DP_OP_20J1_122_6644_n117 n365 A7  n364 FAx1_ASAP7_75t_R
XU508 VSS VDD  n167 n364 N108 NOR2xp33_ASAP7_75t_R
XU509 VSS VDD  n190 DP_OP_20J1_122_6644_n117 DP_OP_20J1_122_6644_n114 n368 MAJIxp5_ASAP7_75t_R
XU510 VSS VDD  DP_OP_20J1_122_6644_n85 n159 A8  n366 HAxp5_ASAP7_75t_R
XU511 VSS VDD  n368 n366 A9  n367 HAxp5_ASAP7_75t_R
XU512 VSS VDD  n167 n367 N109 NOR2xp33_ASAP7_75t_R
XU513 VSS VDD  n239 DP_OP_20J1_122_6644_n85 n368 n371 MAJIxp5_ASAP7_75t_R
XU514 VSS VDD  DP_OP_20J1_122_6644_n64 n371 n369 XOR2xp5_ASAP7_75t_R
XU515 VSS VDD  n238 n371 DP_OP_20J1_122_6644_n64 n374 MAJIxp5_ASAP7_75t_R
XU516 VSS VDD  DP_OP_20J1_122_6644_n60 n374 n372 XOR2xp5_ASAP7_75t_R
XU517 VSS VDD  DP_OP_20J1_122_6644_n44 n372 A10  n373 HAxp5_ASAP7_75t_R
XU518 VSS VDD  n167 n373 N111 NOR2xp33_ASAP7_75t_R
XU519 VSS VDD  DP_OP_20J1_122_6644_n60 DP_OP_20J1_122_6644_n44 n374 n377 MAJx2_ASAP7_75t_R
XU520 VSS VDD  DP_OP_20J1_122_6644_n43 n377 n375 XOR2xp5_ASAP7_75t_R
XU521 VSS VDD  DP_OP_20J1_122_6644_n39 n375 A11  n376 HAxp5_ASAP7_75t_R
XU522 VSS VDD  n167 n376 N112 NOR2xp33_ASAP7_75t_R
XU523 VSS VDD  DP_OP_20J1_122_6644_n39 DP_OP_20J1_122_6644_n43 n377 n381 MAJIxp5_ASAP7_75t_R
XU524 VSS VDD  DP_OP_20J1_122_6644_n41 n381 n378 XOR2xp5_ASAP7_75t_R
XU525 VSS VDD  n167 n379 N113 NOR2xp33_ASAP7_75t_R
XU526 VSS VDD  n380 DP_OP_20J1_122_6644_n41 n381 n382 MAJIxp5_ASAP7_75t_R
XU527 VSS VDD  n166 n382 N114 AND2x2_ASAP7_75t_R
XU528 VSS VDD  n205 in_valid n384 NOR2xp33_ASAP7_75t_R
XU529 VSS VDD  n204 n384 n150 NOR2xp33_ASAP7_75t_R
XU530 VSS VDD  n166 n386 n149 NOR2xp33_ASAP7_75t_R
.ENDS


