.SUBCKT Convolution_pipeline VSS VDD  clk rst_n in_valid n190 n371 In_IFM_1[3] In_IFM_1[2] In_IFM_1[1] In_IFM_1[0] In_IFM_2[3] In_IFM_2[2] In_IFM_2[1] In_IFM_2[0] In_IFM_3[3] In_IFM_3[2] In_IFM_3[1] In_IFM_3[0] In_IFM_4[3] In_IFM_4[2] In_IFM_4[1] In_IFM_4[0] In_Weight_1[3] In_Weight_1[2] In_Weight_1[1] In_Weight_1[0] In_Weight_2[3] In_Weight_2[2] In_Weight_2[1] In_Weight_2[0] In_Weight_3[3] In_Weight_3[2] In_Weight_3[1] In_Weight_3[0] In_Weight_4[3] In_Weight_4[2] In_Weight_4[1] In_Weight_4[0] Out_OFM[11] Out_OFM[10] Out_OFM[9] Out_OFM[8] Out_OFM[7] Out_OFM[6] Out_OFM[5] Out_OFM[4] Out_OFM[3] Out_OFM[2] Out_OFM[1] Out_OFM[0]
XOut_OFM_reg_9_ VSS VDD  n373 clk n436 n511 n372 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_8_ VSS VDD  n371 clk n436 n557 n370 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_7_ VSS VDD  n369 clk n436 n519 n368 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_6_ VSS VDD  n367 clk n436 n517 n366 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_5_ VSS VDD  n365 clk n436 n484 n364 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_4_ VSS VDD  n363 clk n436 n483 n362 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_3_ VSS VDD  n361 clk n436 n551 n360 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_2_ VSS VDD  n359 clk n436 n523 n358 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_1_ VSS VDD  n357 clk n436 n493 n356 ASYNC_DFFHx1_ASAP7_75t_R
XOut_OFM_reg_0_ VSS VDD  n355 clk n436 n482 n354 ASYNC_DFFHx1_ASAP7_75t_R
XIn_1_reg_3_ VSS VDD  n353 clk n436 n486 n352 ASYNC_DFFHx1_ASAP7_75t_R
XIn_1_reg_2_ VSS VDD  n351 clk n436 n452 n350 ASYNC_DFFHx1_ASAP7_75t_R
XIn_1_reg_1_ VSS VDD  n349 clk n436 n513 n348 ASYNC_DFFHx1_ASAP7_75t_R
XIn_1_reg_0_ VSS VDD  n347 clk n436 n476 n346 ASYNC_DFFHx1_ASAP7_75t_R
XIn_2_reg_3_ VSS VDD  n345 clk n436 n450 n344 ASYNC_DFFHx1_ASAP7_75t_R
XIn_2_reg_2_ VSS VDD  n343 clk n436 n525 n342 ASYNC_DFFHx1_ASAP7_75t_R
XIn_2_reg_1_ VSS VDD  n341 clk n436 n456 n340 ASYNC_DFFHx1_ASAP7_75t_R
XIn_2_reg_0_ VSS VDD  n339 clk n436 n479 n338 ASYNC_DFFHx1_ASAP7_75t_R
XIn_3_reg_3_ VSS VDD  n337 clk n436 n489 n336 ASYNC_DFFHx1_ASAP7_75t_R
XIn_3_reg_2_ VSS VDD  n335 clk n436 n504 n334 ASYNC_DFFHx1_ASAP7_75t_R
XIn_3_reg_1_ VSS VDD  n333 clk n436 n460 n332 ASYNC_DFFHx1_ASAP7_75t_R
XIn_3_reg_0_ VSS VDD  n331 clk n436 n522 n330 ASYNC_DFFHx1_ASAP7_75t_R
XIn_4_reg_3_ VSS VDD  n329 clk n436 n462 n328 ASYNC_DFFHx1_ASAP7_75t_R
XIn_4_reg_2_ VSS VDD  n327 clk n436 n449 n326 ASYNC_DFFHx1_ASAP7_75t_R
XIn_4_reg_1_ VSS VDD  n325 clk n436 n481 n324 ASYNC_DFFHx1_ASAP7_75t_R
XIn_4_reg_0_ VSS VDD  n323 clk n436 n453 n322 ASYNC_DFFHx1_ASAP7_75t_R
Xweight1_reg_3_ VSS VDD  n321 clk n436 n478 n320 ASYNC_DFFHx1_ASAP7_75t_R
Xweight1_reg_2_ VSS VDD  n319 clk n436 n471 n318 ASYNC_DFFHx1_ASAP7_75t_R
Xweight1_reg_1_ VSS VDD  n317 clk n436 n495 n316 ASYNC_DFFHx1_ASAP7_75t_R
Xweight1_reg_0_ VSS VDD  n315 clk n436 n464 n314 ASYNC_DFFHx1_ASAP7_75t_R
Xweight2_reg_3_ VSS VDD  n313 clk n436 n524 n312 ASYNC_DFFHx1_ASAP7_75t_R
Xweight2_reg_2_ VSS VDD  n311 clk n436 n488 n310 ASYNC_DFFHx1_ASAP7_75t_R
Xweight2_reg_1_ VSS VDD  n309 clk n436 n558 n308 ASYNC_DFFHx1_ASAP7_75t_R
Xweight2_reg_0_ VSS VDD  n307 clk n436 n463 n306 ASYNC_DFFHx1_ASAP7_75t_R
Xweight3_reg_3_ VSS VDD  n305 clk n436 n470 n304 ASYNC_DFFHx1_ASAP7_75t_R
Xweight3_reg_2_ VSS VDD  n303 clk n436 n499 n302 ASYNC_DFFHx1_ASAP7_75t_R
Xweight3_reg_1_ VSS VDD  n301 clk n436 n487 n300 ASYNC_DFFHx1_ASAP7_75t_R
Xweight3_reg_0_ VSS VDD  n299 clk n436 n506 n298 ASYNC_DFFHx1_ASAP7_75t_R
Xweight4_reg_3_ VSS VDD  n297 clk n436 n468 n296 ASYNC_DFFHx1_ASAP7_75t_R
Xweight4_reg_2_ VSS VDD  n295 clk n436 n490 n294 ASYNC_DFFHx1_ASAP7_75t_R
Xweight4_reg_1_ VSS VDD  n293 clk n436 n451 n292 ASYNC_DFFHx1_ASAP7_75t_R
Xweight4_reg_0_ VSS VDD  n291 clk n436 n466 n290 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_1_reg_7_ VSS VDD  n289 clk n436 n516 n288 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_1_reg_6_ VSS VDD  n287 clk n436 n510 n286 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_1_reg_5_ VSS VDD  n285 clk n436 n553 n284 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_1_reg_4_ VSS VDD  n283 clk n436 n528 n282 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_1_reg_3_ VSS VDD  n281 clk n436 n515 n280 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_1_reg_2_ VSS VDD  n279 clk n436 n526 n278 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_1_reg_1_ VSS VDD  n277 clk n436 n552 n276 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_1_reg_0_ VSS VDD  n275 clk n436 n512 n274 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_2_reg_7_ VSS VDD  n273 clk n436 n500 n272 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_2_reg_6_ VSS VDD  n271 clk n436 n494 n270 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_2_reg_5_ VSS VDD  n269 clk n436 n448 n268 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_2_reg_4_ VSS VDD  n267 clk n436 n518 n266 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_2_reg_3_ VSS VDD  n265 clk n436 n507 n264 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_2_reg_2_ VSS VDD  n263 clk n436 n492 n262 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_2_reg_1_ VSS VDD  n261 clk n436 n480 n260 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_2_reg_0_ VSS VDD  n259 clk n436 n501 n258 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_3_reg_7_ VSS VDD  n257 clk n436 n527 n256 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_3_reg_6_ VSS VDD  n255 clk n436 n458 n254 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_3_reg_5_ VSS VDD  n253 clk n436 n542 n252 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_3_reg_4_ VSS VDD  n251 clk n436 n467 n250 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_3_reg_3_ VSS VDD  n249 clk n436 n455 n248 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_3_reg_2_ VSS VDD  n247 clk n436 n521 n246 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_3_reg_1_ VSS VDD  n245 clk n436 n469 n244 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_3_reg_0_ VSS VDD  n243 clk n436 n475 n242 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_4_reg_7_ VSS VDD  n241 clk n436 n491 n240 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_4_reg_6_ VSS VDD  n239 clk n436 n529 n238 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_4_reg_5_ VSS VDD  n237 clk n436 n496 n236 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_4_reg_4_ VSS VDD  n235 clk n436 n505 n234 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_4_reg_3_ VSS VDD  n233 clk n436 n457 n232 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_4_reg_2_ VSS VDD  n231 clk n436 n559 n230 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_4_reg_1_ VSS VDD  n229 clk n436 n465 n228 ASYNC_DFFHx1_ASAP7_75t_R
XPPR1_4_reg_0_ VSS VDD  n227 clk n436 n497 n226 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_1_reg_8_ VSS VDD  n225 clk n436 n536 n224 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_1_reg_7_ VSS VDD  n223 clk n436 n477 n222 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_1_reg_6_ VSS VDD  n221 clk n436 n520 n220 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_1_reg_5_ VSS VDD  n219 clk n436 n514 n218 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_1_reg_4_ VSS VDD  n217 clk n436 n556 n216 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_1_reg_3_ VSS VDD  n215 clk n436 n535 n214 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_1_reg_2_ VSS VDD  n213 clk n436 n461 n212 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_1_reg_1_ VSS VDD  n211 clk n436 n498 n210 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_1_reg_0_ VSS VDD  n209 clk n436 n472 n208 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_2_reg_8_ VSS VDD  n207 clk n436 n543 n206 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_2_reg_7_ VSS VDD  n205 clk n436 n554 n204 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_2_reg_6_ VSS VDD  n203 clk n436 n473 n202 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_2_reg_5_ VSS VDD  n201 clk n436 n485 n200 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_2_reg_4_ VSS VDD  n199 clk n436 n502 n198 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_2_reg_3_ VSS VDD  n197 clk n436 n459 n196 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_2_reg_2_ VSS VDD  n195 clk n436 n503 n194 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_2_reg_1_ VSS VDD  n193 clk n436 n474 n192 ASYNC_DFFHx1_ASAP7_75t_R
XPPR2_2_reg_0_ VSS VDD  n191 clk n436 n454 n190 ASYNC_DFFHx1_ASAP7_75t_R
Xmult_x_4_U39 VSS VDD  mult_x_4_n49 mult_x_4_n52 mult_x_4_n38 mult_x_4_n34 mult_x_4_n35 FAx1_ASAP7_75t_R
Xmult_x_4_U35 VSS VDD  mult_x_4_n36 mult_x_4_n45 mult_x_4_n32 mult_x_4_n29 mult_x_4_n30 FAx1_ASAP7_75t_R
Xmult_x_4_U32 VSS VDD  mult_x_4_n41 mult_x_4_n44 mult_x_4_n31 mult_x_4_n25 mult_x_4_n26 FAx1_ASAP7_75t_R
Xmult_x_3_U39 VSS VDD  mult_x_3_n49 mult_x_3_n52 mult_x_3_n38 mult_x_3_n34 mult_x_3_n35 FAx1_ASAP7_75t_R
Xmult_x_3_U35 VSS VDD  mult_x_3_n36 mult_x_3_n45 mult_x_3_n32 mult_x_3_n29 mult_x_3_n30 FAx1_ASAP7_75t_R
Xmult_x_3_U32 VSS VDD  mult_x_3_n41 mult_x_3_n44 mult_x_3_n31 mult_x_3_n25 mult_x_3_n26 FAx1_ASAP7_75t_R
Xmult_x_2_U39 VSS VDD  mult_x_2_n49 mult_x_2_n52 mult_x_2_n38 mult_x_2_n34 mult_x_2_n35 FAx1_ASAP7_75t_R
Xmult_x_2_U35 VSS VDD  mult_x_2_n36 mult_x_2_n45 mult_x_2_n32 mult_x_2_n29 mult_x_2_n30 FAx1_ASAP7_75t_R
Xmult_x_2_U32 VSS VDD  mult_x_2_n41 mult_x_2_n44 mult_x_2_n31 mult_x_2_n25 mult_x_2_n26 FAx1_ASAP7_75t_R
Xmult_x_1_U39 VSS VDD  mult_x_1_n49 mult_x_1_n52 mult_x_1_n38 mult_x_1_n34 mult_x_1_n35 FAx1_ASAP7_75t_R
Xmult_x_1_U35 VSS VDD  mult_x_1_n36 mult_x_1_n45 mult_x_1_n32 mult_x_1_n29 mult_x_1_n30 FAx1_ASAP7_75t_R
Xmult_x_1_U32 VSS VDD  mult_x_1_n41 mult_x_1_n44 mult_x_1_n31 mult_x_1_n25 mult_x_1_n26 FAx1_ASAP7_75t_R
XU381 VSS VDD  n974 n973 n975 NOR2xp33_ASAP7_75t_R
XU382 VSS VDD  n546 n545 INVx2_ASAP7_75t_R
XU383 VSS VDD  n587 n936 INVx2_ASAP7_75t_R
XU384 VSS VDD  n586 n931 INVx2_ASAP7_75t_R
XU385 VSS VDD  n588 n926 INVx2_ASAP7_75t_R
XU386 VSS VDD  n585 n942 INVx2_ASAP7_75t_R
XU387 VSS VDD  mult_x_2_n36 n813 n867 NOR2xp33_ASAP7_75t_R
XU388 VSS VDD  mult_x_4_n36 n791 n857 NOR2xp33_ASAP7_75t_R
XU389 VSS VDD  mult_x_1_n36 n802 n862 NOR2xp33_ASAP7_75t_R
XU390 VSS VDD  n539 n538 INVx2_ASAP7_75t_R
XU391 VSS VDD  n550 n549 INVx2_ASAP7_75t_R
XU392 VSS VDD  n541 n540 INVx2_ASAP7_75t_R
XU393 VSS VDD  n548 n547 INVx2_ASAP7_75t_R
XU394 VSS VDD  n344 n586 BUFx5_ASAP7_75t_R
XU395 VSS VDD  n336 n587 BUFx5_ASAP7_75t_R
XU396 VSS VDD  n328 n588 BUFx5_ASAP7_75t_R
XU397 VSS VDD  n352 n585 BUFx5_ASAP7_75t_R
XU398 VSS VDD  n258 n274 n704 NOR2xp33_ASAP7_75t_R
XU399 VSS VDD  n226 n242 n711 NOR2xp33_ASAP7_75t_R
XU400 VSS VDD  n190 n208 n718 NOR2xp33_ASAP7_75t_R
XU401 VSS VDD  n350 n428 BUFx5_ASAP7_75t_R
XU402 VSS VDD  n326 n425 BUFx5_ASAP7_75t_R
XU403 VSS VDD  n304 n426 BUFx5_ASAP7_75t_R
XU404 VSS VDD  n296 n430 BUFx5_ASAP7_75t_R
XU405 VSS VDD  n342 n429 BUFx5_ASAP7_75t_R
XU406 VSS VDD  n334 n427 BUFx5_ASAP7_75t_R
XU407 VSS VDD  n320 n431 BUFx5_ASAP7_75t_R
XU408 VSS VDD  n582 n421 INVx3_ASAP7_75t_R
XU409 VSS VDD  n581 n422 INVx3_ASAP7_75t_R
XU410 VSS VDD  n584 n423 INVx3_ASAP7_75t_R
XU411 VSS VDD  n583 n424 INVx3_ASAP7_75t_R
XU412 VSS VDD  n256 n580 BUFx5_ASAP7_75t_R
XU413 VSS VDD  n288 n579 BUFx5_ASAP7_75t_R
XU414 VSS VDD  in_valid n379 INVx8_ASAP7_75t_R
XU415 VSS VDD  in_valid n380 INVx8_ASAP7_75t_R
XU416 VSS VDD  in_valid n381 INVx8_ASAP7_75t_R
XU417 VSS VDD  in_valid n382 INVx8_ASAP7_75t_R
XU418 VSS VDD  in_valid n383 INVx8_ASAP7_75t_R
XU419 VSS VDD  in_valid n384 INVx8_ASAP7_75t_R
XU420 VSS VDD  in_valid n385 INVx8_ASAP7_75t_R
XU421 VSS VDD  in_valid n386 INVx8_ASAP7_75t_R
XU422 VSS VDD  in_valid n387 INVx8_ASAP7_75t_R
XU423 VSS VDD  in_valid n388 INVx8_ASAP7_75t_R
XU424 VSS VDD  in_valid n389 INVx8_ASAP7_75t_R
XU425 VSS VDD  in_valid n390 INVx8_ASAP7_75t_R
XU426 VSS VDD  in_valid n391 INVx8_ASAP7_75t_R
XU427 VSS VDD  in_valid n392 INVx8_ASAP7_75t_R
XU428 VSS VDD  in_valid n393 INVx8_ASAP7_75t_R
XU429 VSS VDD  in_valid n394 INVx8_ASAP7_75t_R
XU430 VSS VDD  in_valid n395 INVx8_ASAP7_75t_R
XU431 VSS VDD  in_valid n396 INVx8_ASAP7_75t_R
XU432 VSS VDD  in_valid n397 INVx8_ASAP7_75t_R
XU433 VSS VDD  in_valid n398 INVx8_ASAP7_75t_R
XU434 VSS VDD  in_valid n399 INVx8_ASAP7_75t_R
XU435 VSS VDD  in_valid n400 INVx8_ASAP7_75t_R
XU436 VSS VDD  in_valid n401 INVx8_ASAP7_75t_R
XU437 VSS VDD  in_valid n402 INVx8_ASAP7_75t_R
XU438 VSS VDD  in_valid n403 INVx8_ASAP7_75t_R
XU439 VSS VDD  in_valid n404 INVx8_ASAP7_75t_R
XU440 VSS VDD  in_valid n405 INVx8_ASAP7_75t_R
XU441 VSS VDD  in_valid n406 INVx8_ASAP7_75t_R
XU442 VSS VDD  in_valid n407 INVx8_ASAP7_75t_R
XU443 VSS VDD  in_valid n408 INVx8_ASAP7_75t_R
XU444 VSS VDD  in_valid n409 INVx8_ASAP7_75t_R
XU445 VSS VDD  in_valid n410 INVx8_ASAP7_75t_R
XU446 VSS VDD  in_valid n411 INVx8_ASAP7_75t_R
XU447 VSS VDD  in_valid n412 INVx8_ASAP7_75t_R
XU448 VSS VDD  in_valid n413 INVx8_ASAP7_75t_R
XU449 VSS VDD  in_valid n414 INVx8_ASAP7_75t_R
XU450 VSS VDD  in_valid n415 INVx8_ASAP7_75t_R
XU451 VSS VDD  in_valid n416 INVx8_ASAP7_75t_R
XU452 VSS VDD  in_valid n417 INVx8_ASAP7_75t_R
XU453 VSS VDD  in_valid n418 INVx8_ASAP7_75t_R
XU454 VSS VDD  mult_x_3_n35 n583 BUFx4_ASAP7_75t_R
XU455 VSS VDD  n924 n923 n373 NAND2xp33_ASAP7_75t_R
XU456 VSS VDD  mult_x_2_n35 n582 BUFx4_ASAP7_75t_R
XU457 VSS VDD  mult_x_1_n35 n581 BUFx4_ASAP7_75t_R
XU458 VSS VDD  mult_x_4_n35 n584 BUFx4_ASAP7_75t_R
XU459 VSS VDD  n875 n874 n365 NAND2xp33_ASAP7_75t_R
XU460 VSS VDD  n894 n893 n367 NAND2xp33_ASAP7_75t_R
XU461 VSS VDD  n951 n950 n369 NAND2xp33_ASAP7_75t_R
XU462 VSS VDD  n978 n977 n371 NAND2xp33_ASAP7_75t_R
XU463 VSS VDD  n701 n700 n357 NAND2xp33_ASAP7_75t_R
XU464 VSS VDD  n722 n721 n359 NAND2xp33_ASAP7_75t_R
XU465 VSS VDD  n778 n777 n363 NAND2xp33_ASAP7_75t_R
XU466 VSS VDD  n692 n691 n355 NAND2xp33_ASAP7_75t_R
XU467 VSS VDD  n639 n638 n353 NAND2xp33_ASAP7_75t_R
XU468 VSS VDD  n637 n636 n337 NAND2xp33_ASAP7_75t_R
XU469 VSS VDD  n593 n592 n343 NAND2xp33_ASAP7_75t_R
XU470 VSS VDD  n633 n632 n345 NAND2xp33_ASAP7_75t_R
XU471 VSS VDD  n595 n594 n351 NAND2xp33_ASAP7_75t_R
XU472 VSS VDD  n615 n614 n321 NAND2xp33_ASAP7_75t_R
XU473 VSS VDD  n597 n596 n327 NAND2xp33_ASAP7_75t_R
XU474 VSS VDD  n635 n634 n329 NAND2xp33_ASAP7_75t_R
XU475 VSS VDD  n599 n598 n335 NAND2xp33_ASAP7_75t_R
XU476 VSS VDD  n607 n606 n305 NAND2xp33_ASAP7_75t_R
XU477 VSS VDD  n611 n610 n307 NAND2xp33_ASAP7_75t_R
XU478 VSS VDD  n605 n604 n313 NAND2xp33_ASAP7_75t_R
XU479 VSS VDD  n613 n612 n315 NAND2xp33_ASAP7_75t_R
XU480 VSS VDD  n900 n899 n285 NAND2xp33_ASAP7_75t_R
XU481 VSS VDD  n603 n602 n291 NAND2xp33_ASAP7_75t_R
XU482 VSS VDD  n601 n600 n297 NAND2xp33_ASAP7_75t_R
XU483 VSS VDD  n609 n608 n299 NAND2xp33_ASAP7_75t_R
XU484 VSS VDD  n821 n820 n265 NAND2xp33_ASAP7_75t_R
XU485 VSS VDD  n912 n911 n269 NAND2xp33_ASAP7_75t_R
XU486 VSS VDD  n679 n678 n277 NAND2xp33_ASAP7_75t_R
XU487 VSS VDD  n810 n809 n281 NAND2xp33_ASAP7_75t_R
XU488 VSS VDD  n689 n688 n245 NAND2xp33_ASAP7_75t_R
XU489 VSS VDD  n832 n831 n249 NAND2xp33_ASAP7_75t_R
XU490 VSS VDD  n906 n905 n253 NAND2xp33_ASAP7_75t_R
XU491 VSS VDD  n684 n683 n261 NAND2xp33_ASAP7_75t_R
XU492 VSS VDD  n881 n880 n223 NAND2xp33_ASAP7_75t_R
XU493 VSS VDD  n674 n673 n229 NAND2xp33_ASAP7_75t_R
XU494 VSS VDD  n799 n798 n233 NAND2xp33_ASAP7_75t_R
XU495 VSS VDD  n918 n917 n237 NAND2xp33_ASAP7_75t_R
XU496 VSS VDD  n887 n886 n205 NAND2xp33_ASAP7_75t_R
XU497 VSS VDD  n727 n726 n215 NAND2xp33_ASAP7_75t_R
XU498 VSS VDD  n788 n787 n219 NAND2xp33_ASAP7_75t_R
XU499 VSS VDD  n698 n697 n193 NAND2xp33_ASAP7_75t_R
XU500 VSS VDD  n732 n731 n197 NAND2xp33_ASAP7_75t_R
XU501 VSS VDD  n783 n782 n201 NAND2xp33_ASAP7_75t_R
XU502 VSS VDD  n940 n939 n257 NAND2xp33_ASAP7_75t_R
XU503 VSS VDD  n946 n945 n289 NAND2xp33_ASAP7_75t_R
XU504 VSS VDD  in_valid n419 INVx8_ASAP7_75t_R
XU505 VSS VDD  in_valid n420 INVx8_ASAP7_75t_R
XU506 VSS VDD  n306 n539 BUFx5_ASAP7_75t_R
XU507 VSS VDD  n298 n550 BUFx5_ASAP7_75t_R
XU508 VSS VDD  n312 n546 BUFx5_ASAP7_75t_R
XU509 VSS VDD  n314 n541 BUFx5_ASAP7_75t_R
XU510 VSS VDD  n290 n548 BUFx5_ASAP7_75t_R
XU511 VSS VDD  in_valid n432 INVx8_ASAP7_75t_R
XU512 VSS VDD  in_valid n433 INVx8_ASAP7_75t_R
XU513 VSS VDD  in_valid n434 INVx8_ASAP7_75t_R
XU514 VSS VDD  in_valid n435 INVx8_ASAP7_75t_R
XU515 VSS VDD  in_valid n441 INVx8_ASAP7_75t_R
XU516 VSS VDD  in_valid n440 INVx8_ASAP7_75t_R
XU517 VSS VDD  mult_x_3_n36 n824 n852 NOR2xp33_ASAP7_75t_R
XU518 VSS VDD  n735 n734 n803 NAND2xp33_ASAP7_75t_R
XU519 VSS VDD  n695 n694 n211 NAND2xp33_ASAP7_75t_R
XU520 VSS VDD  n929 n928 n241 NAND2xp33_ASAP7_75t_R
XU521 VSS VDD  n971 n970 n271 NAND2xp33_ASAP7_75t_R
XU522 VSS VDD  n653 n652 n301 NAND2xp33_ASAP7_75t_R
XU523 VSS VDD  n617 n616 n331 NAND2xp33_ASAP7_75t_R
XU524 VSS VDD  n761 n760 n361 NAND2xp33_ASAP7_75t_R
XU525 VSS VDD  n354 Out_OFM[0] INVxp67_ASAP7_75t_R
XU526 VSS VDD  n372 Out_OFM[9] INVxp67_ASAP7_75t_R
XU527 VSS VDD  n368 Out_OFM[7] INVxp67_ASAP7_75t_R
XU528 VSS VDD  n956 n955 n255 NAND2xp5_ASAP7_75t_R
XU529 VSS VDD  n961 n960 n239 NAND2xp5_ASAP7_75t_R
XU530 VSS VDD  n966 n965 n287 NAND2xp5_ASAP7_75t_R
XU531 VSS VDD  n934 n933 n273 NAND2xp5_ASAP7_75t_R
XU532 VSS VDD  n850 n849 n203 NAND2xp5_ASAP7_75t_R
XU533 VSS VDD  n845 n844 n221 NAND2xp5_ASAP7_75t_R
XU534 VSS VDD  n836 n835 n207 NAND2xp5_ASAP7_75t_R
XU535 VSS VDD  n860 n859 n235 NAND2xp5_ASAP7_75t_R
XU536 VSS VDD  n855 n854 n251 NAND2xp5_ASAP7_75t_R
XU537 VSS VDD  n840 n839 n225 NAND2xp5_ASAP7_75t_R
XU538 VSS VDD  n865 n864 n283 NAND2xp5_ASAP7_75t_R
XU539 VSS VDD  n870 n869 n267 NAND2xp5_ASAP7_75t_R
XU540 VSS VDD  n877 n876 n878 NAND2xp5_ASAP7_75t_R
XU541 VSS VDD  n883 n882 n884 NAND2xp5_ASAP7_75t_R
XU542 VSS VDD  n771 n770 n217 NAND2xp5_ASAP7_75t_R
XU543 VSS VDD  n766 n765 n199 NAND2xp5_ASAP7_75t_R
XU544 VSS VDD  n738 n737 n279 NAND2xp5_ASAP7_75t_R
XU545 VSS VDD  n750 n749 n247 NAND2xp5_ASAP7_75t_R
XU546 VSS VDD  n756 n755 n263 NAND2xp5_ASAP7_75t_R
XU547 VSS VDD  n715 n714 n195 NAND2xp5_ASAP7_75t_R
XU548 VSS VDD  n744 n743 n231 NAND2xp5_ASAP7_75t_R
XU549 VSS VDD  n708 n707 n213 NAND2xp5_ASAP7_75t_R
XU550 VSS VDD  n663 n662 n275 NAND2xp5_ASAP7_75t_R
XU551 VSS VDD  n661 n660 n243 NAND2xp5_ASAP7_75t_R
XU552 VSS VDD  n659 n658 n227 NAND2xp5_ASAP7_75t_R
XU553 VSS VDD  n657 n656 n259 NAND2xp5_ASAP7_75t_R
XU554 VSS VDD  n753 n752 n814 NAND2xp5_ASAP7_75t_R
XU555 VSS VDD  n747 n746 n825 NAND2xp5_ASAP7_75t_R
XU556 VSS VDD  n741 n740 n792 NAND2xp5_ASAP7_75t_R
XU557 VSS VDD  n426 n561 INVx2_ASAP7_75t_R
XU558 VSS VDD  n666 n665 n209 NAND2xp5_ASAP7_75t_R
XU559 VSS VDD  n430 n560 INVx2_ASAP7_75t_R
XU560 VSS VDD  n431 n562 INVx2_ASAP7_75t_R
XU561 VSS VDD  n669 n668 n191 NAND2xp5_ASAP7_75t_R
XU562 VSS VDD  n651 n650 n309 NAND2xp5_ASAP7_75t_R
XU563 VSS VDD  n619 n618 n339 NAND2xp5_ASAP7_75t_R
XU564 VSS VDD  n641 n640 n341 NAND2xp5_ASAP7_75t_R
XU565 VSS VDD  n631 n630 n295 NAND2xp5_ASAP7_75t_R
XU566 VSS VDD  n625 n624 n311 NAND2xp5_ASAP7_75t_R
XU567 VSS VDD  n627 n626 n303 NAND2xp5_ASAP7_75t_R
XU568 VSS VDD  n655 n654 n293 NAND2xp5_ASAP7_75t_R
XU569 VSS VDD  n649 n648 n317 NAND2xp5_ASAP7_75t_R
XU570 VSS VDD  n629 n628 n319 NAND2xp5_ASAP7_75t_R
XU571 VSS VDD  n645 n644 n333 NAND2xp5_ASAP7_75t_R
XU572 VSS VDD  n623 n622 n323 NAND2xp5_ASAP7_75t_R
XU573 VSS VDD  n647 n646 n325 NAND2xp5_ASAP7_75t_R
XU574 VSS VDD  n621 n620 n347 NAND2xp5_ASAP7_75t_R
XU575 VSS VDD  n643 n642 n349 NAND2xp5_ASAP7_75t_R
XU576 VSS VDD  n888 n573 INVx3_ASAP7_75t_R
XU577 VSS VDD  n920 n572 INVx3_ASAP7_75t_R
XU578 VSS VDD  n428 n544 INVx2_ASAP7_75t_R
XU579 VSS VDD  n702 n534 INVx3_ASAP7_75t_R
XU580 VSS VDD  n427 n564 INVx2_ASAP7_75t_R
XU581 VSS VDD  n425 n563 INVx2_ASAP7_75t_R
XU582 VSS VDD  n568 n797 INVx3_ASAP7_75t_R
XU583 VSS VDD  n580 n938 INVx2_ASAP7_75t_R
XU584 VSS VDD  n772 n574 INVx3_ASAP7_75t_R
XU585 VSS VDD  n567 n916 INVx3_ASAP7_75t_R
XU586 VSS VDD  n579 n944 INVx2_ASAP7_75t_R
XU587 VSS VDD  n709 n532 INVx3_ASAP7_75t_R
XU588 VSS VDD  n566 n819 INVx3_ASAP7_75t_R
XU589 VSS VDD  n429 n555 INVx2_ASAP7_75t_R
XU590 VSS VDD  n717 n537 INVx3_ASAP7_75t_R
XU591 VSS VDD  n565 n910 INVx3_ASAP7_75t_R
XU592 VSS VDD  n370 Out_OFM[8] INVxp67_ASAP7_75t_R
XU593 VSS VDD  n360 Out_OFM[3] INVxp67_ASAP7_75t_R
XU594 VSS VDD  n362 Out_OFM[4] INVxp67_ASAP7_75t_R
XU595 VSS VDD  n364 Out_OFM[5] INVxp67_ASAP7_75t_R
XU596 VSS VDD  n358 Out_OFM[2] INVxp67_ASAP7_75t_R
XU597 VSS VDD  n356 Out_OFM[1] INVxp67_ASAP7_75t_R
XU598 VSS VDD  n366 Out_OFM[6] INVxp67_ASAP7_75t_R
XU599 VSS VDD  n436 TIELOx1_ASAP7_75t_R
XU600 VSS VDD  n439 TIEHIx1_ASAP7_75t_R
XU601 VSS VDD  n439 Out_OFM[10] INVxp33_ASAP7_75t_R
XU602 VSS VDD  n439 Out_OFM[11] INVxp33_ASAP7_75t_R
XU603 VSS VDD  n244 n709 BUFx5_ASAP7_75t_R
XU604 VSS VDD  n276 n702 BUFx5_ASAP7_75t_R
XU605 VSS VDD  n210 n717 BUFx5_ASAP7_75t_R
XU606 VSS VDD  mult_x_1_n30 n895 mult_x_1_n34 n442 MAJIxp5_ASAP7_75t_R
XU607 VSS VDD  mult_x_3_n30 n901 mult_x_3_n34 n443 MAJIxp5_ASAP7_75t_R
XU608 VSS VDD  mult_x_2_n30 n907 mult_x_2_n34 n444 MAJIxp5_ASAP7_75t_R
XU609 VSS VDD  mult_x_4_n30 n913 mult_x_4_n34 n445 MAJIxp5_ASAP7_75t_R
XU610 VSS VDD  mult_x_1_n30 n895 mult_x_1_n34 n941 MAJx2_ASAP7_75t_R
XU611 VSS VDD  mult_x_2_n30 n907 mult_x_2_n34 n930 MAJx2_ASAP7_75t_R
XU612 VSS VDD  mult_x_4_n30 n913 mult_x_4_n34 n925 MAJx2_ASAP7_75t_R
XU613 VSS VDD  mult_x_3_n30 n901 mult_x_3_n34 n935 MAJx2_ASAP7_75t_R
XU614 VSS VDD  n846 n254 n238 n446 MAJIxp5_ASAP7_75t_R
XU615 VSS VDD  n841 n286 n270 n447 MAJIxp5_ASAP7_75t_R
XU616 VSS VDD  rst_n n448 INVx8_ASAP7_75t_R
XU617 VSS VDD  rst_n n449 INVx8_ASAP7_75t_R
XU618 VSS VDD  rst_n n450 INVx8_ASAP7_75t_R
XU619 VSS VDD  rst_n n451 INVx8_ASAP7_75t_R
XU620 VSS VDD  rst_n n452 INVx8_ASAP7_75t_R
XU621 VSS VDD  rst_n n453 INVx8_ASAP7_75t_R
XU622 VSS VDD  rst_n n454 INVx8_ASAP7_75t_R
XU623 VSS VDD  rst_n n455 INVx8_ASAP7_75t_R
XU624 VSS VDD  rst_n n456 INVx8_ASAP7_75t_R
XU625 VSS VDD  rst_n n457 INVx8_ASAP7_75t_R
XU626 VSS VDD  rst_n n458 INVx8_ASAP7_75t_R
XU627 VSS VDD  rst_n n459 INVx8_ASAP7_75t_R
XU628 VSS VDD  rst_n n460 INVx8_ASAP7_75t_R
XU629 VSS VDD  rst_n n461 INVx8_ASAP7_75t_R
XU630 VSS VDD  rst_n n462 INVx8_ASAP7_75t_R
XU631 VSS VDD  rst_n n463 INVx8_ASAP7_75t_R
XU632 VSS VDD  rst_n n464 INVx8_ASAP7_75t_R
XU633 VSS VDD  rst_n n465 INVx8_ASAP7_75t_R
XU634 VSS VDD  rst_n n466 INVx8_ASAP7_75t_R
XU635 VSS VDD  rst_n n467 INVx8_ASAP7_75t_R
XU636 VSS VDD  rst_n n468 INVx8_ASAP7_75t_R
XU637 VSS VDD  rst_n n469 INVx8_ASAP7_75t_R
XU638 VSS VDD  rst_n n470 INVx8_ASAP7_75t_R
XU639 VSS VDD  rst_n n471 INVx8_ASAP7_75t_R
XU640 VSS VDD  rst_n n472 INVx8_ASAP7_75t_R
XU641 VSS VDD  rst_n n473 INVx8_ASAP7_75t_R
XU642 VSS VDD  rst_n n474 INVx8_ASAP7_75t_R
XU643 VSS VDD  rst_n n475 INVx8_ASAP7_75t_R
XU644 VSS VDD  rst_n n476 INVx8_ASAP7_75t_R
XU645 VSS VDD  rst_n n477 INVx8_ASAP7_75t_R
XU646 VSS VDD  rst_n n478 INVx8_ASAP7_75t_R
XU647 VSS VDD  rst_n n479 INVx8_ASAP7_75t_R
XU648 VSS VDD  rst_n n480 INVx8_ASAP7_75t_R
XU649 VSS VDD  rst_n n481 INVx8_ASAP7_75t_R
XU650 VSS VDD  rst_n n482 INVx8_ASAP7_75t_R
XU651 VSS VDD  rst_n n483 INVx8_ASAP7_75t_R
XU652 VSS VDD  rst_n n484 INVx8_ASAP7_75t_R
XU653 VSS VDD  rst_n n485 INVx8_ASAP7_75t_R
XU654 VSS VDD  rst_n n486 INVx8_ASAP7_75t_R
XU655 VSS VDD  rst_n n487 INVx8_ASAP7_75t_R
XU656 VSS VDD  rst_n n488 INVx8_ASAP7_75t_R
XU657 VSS VDD  rst_n n489 INVx8_ASAP7_75t_R
XU658 VSS VDD  rst_n n490 INVx8_ASAP7_75t_R
XU659 VSS VDD  rst_n n491 INVx8_ASAP7_75t_R
XU660 VSS VDD  rst_n n492 INVx8_ASAP7_75t_R
XU661 VSS VDD  rst_n n493 INVx8_ASAP7_75t_R
XU662 VSS VDD  rst_n n494 INVx8_ASAP7_75t_R
XU663 VSS VDD  rst_n n495 INVx8_ASAP7_75t_R
XU664 VSS VDD  rst_n n496 INVx8_ASAP7_75t_R
XU665 VSS VDD  rst_n n497 INVx8_ASAP7_75t_R
XU666 VSS VDD  rst_n n498 INVx8_ASAP7_75t_R
XU667 VSS VDD  rst_n n499 INVx8_ASAP7_75t_R
XU668 VSS VDD  n258 n274 n530 OR2x2_ASAP7_75t_R
XU669 VSS VDD  n226 n242 n531 OR2x2_ASAP7_75t_R
XU670 VSS VDD  n190 n208 n533 OR2x2_ASAP7_75t_R
XU671 VSS VDD  rst_n n500 INVx8_ASAP7_75t_R
XU672 VSS VDD  rst_n n501 INVx8_ASAP7_75t_R
XU673 VSS VDD  rst_n n502 INVx8_ASAP7_75t_R
XU674 VSS VDD  rst_n n503 INVx8_ASAP7_75t_R
XU675 VSS VDD  rst_n n504 INVx8_ASAP7_75t_R
XU676 VSS VDD  rst_n n505 INVx8_ASAP7_75t_R
XU677 VSS VDD  rst_n n506 INVx8_ASAP7_75t_R
XU678 VSS VDD  rst_n n507 INVx8_ASAP7_75t_R
XU679 VSS VDD  n830 n578 INVx3_ASAP7_75t_R
XU680 VSS VDD  n808 n576 INVx3_ASAP7_75t_R
XU681 VSS VDD  n904 n577 INVx3_ASAP7_75t_R
XU682 VSS VDD  n898 n575 INVx3_ASAP7_75t_R
XU683 VSS VDD  n729 n568 n730 XNOR2xp5_ASAP7_75t_R
XU684 VSS VDD  n232 n568 BUFx5_ASAP7_75t_R
XU685 VSS VDD  n222 n569 BUFx5_ASAP7_75t_R
XU686 VSS VDD  n218 n570 BUFx5_ASAP7_75t_R
XU687 VSS VDD  n214 n571 BUFx5_ASAP7_75t_R
XU688 VSS VDD  n724 n566 n725 XNOR2xp5_ASAP7_75t_R
XU689 VSS VDD  n264 n566 BUFx5_ASAP7_75t_R
XU690 VSS VDD  n780 n567 n781 XNOR2xp5_ASAP7_75t_R
XU691 VSS VDD  n236 n567 BUFx5_ASAP7_75t_R
XU692 VSS VDD  n785 n565 n786 XNOR2xp5_ASAP7_75t_R
XU693 VSS VDD  n268 n565 BUFx5_ASAP7_75t_R
XU694 VSS VDD  n846 n254 n238 n508 MAJx2_ASAP7_75t_R
XU695 VSS VDD  n841 n286 n270 n509 MAJx2_ASAP7_75t_R
XU696 VSS VDD  rst_n n510 INVx8_ASAP7_75t_R
XU697 VSS VDD  rst_n n511 INVx8_ASAP7_75t_R
XU698 VSS VDD  rst_n n512 INVx8_ASAP7_75t_R
XU699 VSS VDD  rst_n n513 INVx8_ASAP7_75t_R
XU700 VSS VDD  rst_n n514 INVx8_ASAP7_75t_R
XU701 VSS VDD  rst_n n515 INVx8_ASAP7_75t_R
XU702 VSS VDD  rst_n n516 INVx8_ASAP7_75t_R
XU703 VSS VDD  rst_n n517 INVx8_ASAP7_75t_R
XU704 VSS VDD  rst_n n518 INVx8_ASAP7_75t_R
XU705 VSS VDD  rst_n n519 INVx8_ASAP7_75t_R
XU706 VSS VDD  rst_n n520 INVx8_ASAP7_75t_R
XU707 VSS VDD  rst_n n521 INVx8_ASAP7_75t_R
XU708 VSS VDD  n703 n590 INVx4_ASAP7_75t_R
XU709 VSS VDD  n260 n703 BUFx5_ASAP7_75t_R
XU710 VSS VDD  n710 n591 INVx4_ASAP7_75t_R
XU711 VSS VDD  n228 n710 BUFx5_ASAP7_75t_R
XU712 VSS VDD  n716 n589 INVx4_ASAP7_75t_R
XU713 VSS VDD  n192 n716 BUFx5_ASAP7_75t_R
XU714 VSS VDD  rst_n n522 INVx8_ASAP7_75t_R
XU715 VSS VDD  rst_n n523 INVx8_ASAP7_75t_R
XU716 VSS VDD  n284 n898 BUFx5_ASAP7_75t_R
XU717 VSS VDD  n204 n920 BUFx5_ASAP7_75t_R
XU718 VSS VDD  n248 n830 BUFx5_ASAP7_75t_R
XU719 VSS VDD  n252 n904 BUFx5_ASAP7_75t_R
XU720 VSS VDD  n280 n808 BUFx5_ASAP7_75t_R
XU721 VSS VDD  rst_n n524 INVx8_ASAP7_75t_R
XU722 VSS VDD  rst_n n525 INVx8_ASAP7_75t_R
XU723 VSS VDD  n196 n772 BUFx5_ASAP7_75t_R
XU724 VSS VDD  n200 n888 BUFx5_ASAP7_75t_R
XU725 VSS VDD  rst_n n526 INVx8_ASAP7_75t_R
XU726 VSS VDD  rst_n n527 INVx8_ASAP7_75t_R
XU727 VSS VDD  rst_n n528 INVx8_ASAP7_75t_R
XU728 VSS VDD  rst_n n529 INVx8_ASAP7_75t_R
XU729 VSS VDD  rst_n n535 INVx8_ASAP7_75t_R
XU730 VSS VDD  rst_n n536 INVx8_ASAP7_75t_R
XU731 VSS VDD  rst_n n542 INVx8_ASAP7_75t_R
XU732 VSS VDD  rst_n n543 INVx8_ASAP7_75t_R
XU733 VSS VDD  rst_n n551 INVx8_ASAP7_75t_R
XU734 VSS VDD  rst_n n552 INVx8_ASAP7_75t_R
XU735 VSS VDD  rst_n n553 INVx8_ASAP7_75t_R
XU736 VSS VDD  rst_n n554 INVx8_ASAP7_75t_R
XU737 VSS VDD  rst_n n556 INVx8_ASAP7_75t_R
XU738 VSS VDD  rst_n n557 INVx8_ASAP7_75t_R
XU739 VSS VDD  rst_n n558 INVx8_ASAP7_75t_R
XU740 VSS VDD  rst_n n559 INVx8_ASAP7_75t_R
XU741 VSS VDD  n569 n921 INVx2_ASAP7_75t_R
XU742 VSS VDD  n570 n890 INVx2_ASAP7_75t_R
XU743 VSS VDD  n571 n774 INVx2_ASAP7_75t_R
XU744 VSS VDD  in_valid In_IFM_2[2] n593 NAND2xp33_ASAP7_75t_R
XU745 VSS VDD  n555 n400 n592 NAND2xp33_ASAP7_75t_R
XU746 VSS VDD  in_valid In_IFM_1[2] n595 NAND2xp33_ASAP7_75t_R
XU747 VSS VDD  n544 n379 n594 NAND2xp33_ASAP7_75t_R
XU748 VSS VDD  in_valid In_IFM_4[2] n597 NAND2xp33_ASAP7_75t_R
XU749 VSS VDD  n563 n404 n596 NAND2xp33_ASAP7_75t_R
XU750 VSS VDD  in_valid In_IFM_3[2] n599 NAND2xp33_ASAP7_75t_R
XU751 VSS VDD  n564 n411 n598 NAND2xp33_ASAP7_75t_R
XU752 VSS VDD  in_valid In_Weight_4[3] n601 NAND2xp33_ASAP7_75t_R
XU753 VSS VDD  n560 n434 n600 NAND2xp33_ASAP7_75t_R
XU754 VSS VDD  in_valid In_Weight_4[0] n603 NAND2xp33_ASAP7_75t_R
XU755 VSS VDD  n547 n412 n602 NAND2xp33_ASAP7_75t_R
XU756 VSS VDD  in_valid In_Weight_2[3] n605 NAND2xp33_ASAP7_75t_R
XU757 VSS VDD  n545 n413 n604 NAND2xp33_ASAP7_75t_R
XU758 VSS VDD  in_valid In_Weight_3[3] n607 NAND2xp33_ASAP7_75t_R
XU759 VSS VDD  n561 n399 n606 NAND2xp33_ASAP7_75t_R
XU760 VSS VDD  in_valid In_Weight_3[0] n609 NAND2xp33_ASAP7_75t_R
XU761 VSS VDD  n549 n387 n608 NAND2xp33_ASAP7_75t_R
XU762 VSS VDD  in_valid In_Weight_2[0] n611 NAND2xp33_ASAP7_75t_R
XU763 VSS VDD  n538 n389 n610 NAND2xp33_ASAP7_75t_R
XU764 VSS VDD  in_valid In_Weight_1[0] n613 NAND2xp33_ASAP7_75t_R
XU765 VSS VDD  n540 n397 n612 NAND2xp33_ASAP7_75t_R
XU766 VSS VDD  in_valid In_Weight_1[3] n615 NAND2xp33_ASAP7_75t_R
XU767 VSS VDD  n562 n409 n614 NAND2xp33_ASAP7_75t_R
XU768 VSS VDD  in_valid In_IFM_3[0] n617 NAND2xp33_ASAP7_75t_R
XU769 VSS VDD  in_valid n330 n616 OR2x2_ASAP7_75t_R
XU770 VSS VDD  in_valid In_IFM_2[0] n619 NAND2xp33_ASAP7_75t_R
XU771 VSS VDD  in_valid n338 n618 OR2x2_ASAP7_75t_R
XU772 VSS VDD  in_valid In_IFM_1[0] n621 NAND2xp33_ASAP7_75t_R
XU773 VSS VDD  in_valid n346 n620 OR2x2_ASAP7_75t_R
XU774 VSS VDD  in_valid In_IFM_4[0] n623 NAND2xp33_ASAP7_75t_R
XU775 VSS VDD  in_valid n322 n622 OR2x2_ASAP7_75t_R
XU776 VSS VDD  in_valid In_Weight_2[2] n625 NAND2xp33_ASAP7_75t_R
XU777 VSS VDD  in_valid n310 n624 OR2x2_ASAP7_75t_R
XU778 VSS VDD  in_valid In_Weight_3[2] n627 NAND2xp33_ASAP7_75t_R
XU779 VSS VDD  in_valid n302 n626 OR2x2_ASAP7_75t_R
XU780 VSS VDD  in_valid In_Weight_1[2] n629 NAND2xp33_ASAP7_75t_R
XU781 VSS VDD  in_valid n318 n628 OR2x2_ASAP7_75t_R
XU782 VSS VDD  in_valid In_Weight_4[2] n631 NAND2xp33_ASAP7_75t_R
XU783 VSS VDD  in_valid n294 n630 OR2x2_ASAP7_75t_R
XU784 VSS VDD  in_valid In_IFM_2[3] n633 NAND2xp33_ASAP7_75t_R
XU785 VSS VDD  n931 n386 n632 NAND2xp33_ASAP7_75t_R
XU786 VSS VDD  in_valid In_IFM_4[3] n635 NAND2xp33_ASAP7_75t_R
XU787 VSS VDD  n926 n417 n634 NAND2xp33_ASAP7_75t_R
XU788 VSS VDD  in_valid In_IFM_3[3] n637 NAND2xp33_ASAP7_75t_R
XU789 VSS VDD  n398 n936 n636 NAND2xp33_ASAP7_75t_R
XU790 VSS VDD  in_valid In_IFM_1[3] n639 NAND2xp33_ASAP7_75t_R
XU791 VSS VDD  n942 n396 n638 NAND2xp33_ASAP7_75t_R
XU792 VSS VDD  in_valid In_IFM_2[1] n641 NAND2xp33_ASAP7_75t_R
XU793 VSS VDD  in_valid n340 n640 OR2x2_ASAP7_75t_R
XU794 VSS VDD  in_valid In_IFM_1[1] n643 NAND2xp33_ASAP7_75t_R
XU795 VSS VDD  in_valid n348 n642 OR2x2_ASAP7_75t_R
XU796 VSS VDD  in_valid In_IFM_3[1] n645 NAND2xp33_ASAP7_75t_R
XU797 VSS VDD  in_valid n332 n644 OR2x2_ASAP7_75t_R
XU798 VSS VDD  in_valid In_IFM_4[1] n647 NAND2xp33_ASAP7_75t_R
XU799 VSS VDD  in_valid n324 n646 OR2x2_ASAP7_75t_R
XU800 VSS VDD  in_valid In_Weight_1[1] n649 NAND2xp33_ASAP7_75t_R
XU801 VSS VDD  in_valid n316 n648 OR2x2_ASAP7_75t_R
XU802 VSS VDD  in_valid In_Weight_2[1] n651 NAND2xp33_ASAP7_75t_R
XU803 VSS VDD  in_valid n308 n650 OR2x2_ASAP7_75t_R
XU804 VSS VDD  in_valid In_Weight_3[1] n653 NAND2xp33_ASAP7_75t_R
XU805 VSS VDD  in_valid n300 n652 OR2x2_ASAP7_75t_R
XU806 VSS VDD  in_valid In_Weight_4[1] n655 NAND2xp33_ASAP7_75t_R
XU807 VSS VDD  in_valid n292 n654 OR2x2_ASAP7_75t_R
XU808 VSS VDD  n539 n338 n752 NOR2xp33_ASAP7_75t_R
XU809 VSS VDD  in_valid n752 n657 NAND2xp33_ASAP7_75t_R
XU810 VSS VDD  in_valid n258 n656 OR2x2_ASAP7_75t_R
XU811 VSS VDD  n548 n322 n740 NOR2xp33_ASAP7_75t_R
XU812 VSS VDD  in_valid n740 n659 NAND2xp33_ASAP7_75t_R
XU813 VSS VDD  in_valid n226 n658 OR2x2_ASAP7_75t_R
XU814 VSS VDD  n550 n330 n746 NOR2xp33_ASAP7_75t_R
XU815 VSS VDD  in_valid n746 n661 NAND2xp33_ASAP7_75t_R
XU816 VSS VDD  in_valid n242 n660 OR2x2_ASAP7_75t_R
XU817 VSS VDD  n541 n346 n734 NOR2xp33_ASAP7_75t_R
XU818 VSS VDD  in_valid n734 n663 NAND2xp33_ASAP7_75t_R
XU819 VSS VDD  in_valid n274 n662 OR2x2_ASAP7_75t_R
XU820 VSS VDD  n274 n258 n664 NAND2xp33_ASAP7_75t_R
XU821 VSS VDD  n664 n530 in_valid n666 NAND3xp33_ASAP7_75t_R
XU822 VSS VDD  in_valid n208 n665 OR2x2_ASAP7_75t_R
XU823 VSS VDD  n242 n226 n667 NAND2xp33_ASAP7_75t_R
XU824 VSS VDD  n667 n531 in_valid n669 NAND3xp33_ASAP7_75t_R
XU825 VSS VDD  in_valid n190 n668 OR2x2_ASAP7_75t_R
XU826 VSS VDD  n292 n322 n671 NOR2xp33_ASAP7_75t_R
XU827 VSS VDD  n548 n324 n670 NOR2xp33_ASAP7_75t_R
XU828 VSS VDD  n671 n670 n672 XOR2xp5_ASAP7_75t_R
XU829 VSS VDD  in_valid n672 n674 NAND2xp33_ASAP7_75t_R
XU830 VSS VDD  n591 n380 n673 NAND2xp33_ASAP7_75t_R
XU831 VSS VDD  n316 n346 n676 NOR2xp33_ASAP7_75t_R
XU832 VSS VDD  n541 n348 n675 NOR2xp33_ASAP7_75t_R
XU833 VSS VDD  n676 n675 n677 XOR2xp5_ASAP7_75t_R
XU834 VSS VDD  in_valid n677 n679 NAND2xp33_ASAP7_75t_R
XU835 VSS VDD  n534 n383 n678 NAND2xp33_ASAP7_75t_R
XU836 VSS VDD  n308 n338 n681 NOR2xp33_ASAP7_75t_R
XU837 VSS VDD  n539 n340 n680 NOR2xp33_ASAP7_75t_R
XU838 VSS VDD  n681 n680 n682 XOR2xp5_ASAP7_75t_R
XU839 VSS VDD  in_valid n682 n684 NAND2xp33_ASAP7_75t_R
XU840 VSS VDD  n590 n418 n683 NAND2xp33_ASAP7_75t_R
XU841 VSS VDD  n300 n330 n686 NOR2xp33_ASAP7_75t_R
XU842 VSS VDD  n550 n332 n685 NOR2xp33_ASAP7_75t_R
XU843 VSS VDD  n686 n685 n687 XOR2xp5_ASAP7_75t_R
XU844 VSS VDD  in_valid n687 n689 NAND2xp33_ASAP7_75t_R
XU845 VSS VDD  n532 n384 n688 NAND2xp33_ASAP7_75t_R
XU846 VSS VDD  n208 n190 n690 NAND2xp33_ASAP7_75t_R
XU847 VSS VDD  n690 n533 in_valid n692 NAND3xp33_ASAP7_75t_R
XU848 VSS VDD  Out_OFM[0] n416 n691 NAND2xp33_ASAP7_75t_R
XU849 VSS VDD  n702 n704 n590 A0  n693 FAx1_ASAP7_75t_R
XU850 VSS VDD  in_valid n693 n695 NAND2xp33_ASAP7_75t_R
XU851 VSS VDD  n537 n381 n694 NAND2xp33_ASAP7_75t_R
XU852 VSS VDD  n709 n711 n591 A1  n696 FAx1_ASAP7_75t_R
XU853 VSS VDD  in_valid n696 n698 NAND2xp33_ASAP7_75t_R
XU854 VSS VDD  n589 n385 n697 NAND2xp33_ASAP7_75t_R
XU855 VSS VDD  n717 n718 n589 A2  n699 FAx1_ASAP7_75t_R
XU856 VSS VDD  in_valid n699 n701 NAND2xp33_ASAP7_75t_R
XU857 VSS VDD  Out_OFM[1] n405 n700 NAND2xp33_ASAP7_75t_R
XU858 VSS VDD  n534 n704 n590 n723 MAJIxp5_ASAP7_75t_R
XU859 VSS VDD  n723 n278 n705 XOR2xp5_ASAP7_75t_R
XU860 VSS VDD  n262 n705 A3  n706 HAxp5_ASAP7_75t_R
XU861 VSS VDD  in_valid n706 n708 NAND2xp33_ASAP7_75t_R
XU862 VSS VDD  in_valid n212 n707 OR2x2_ASAP7_75t_R
XU863 VSS VDD  n532 n711 n591 n728 MAJIxp5_ASAP7_75t_R
XU864 VSS VDD  n728 n246 n712 XOR2xp5_ASAP7_75t_R
XU865 VSS VDD  n230 n712 A4  n713 HAxp5_ASAP7_75t_R
XU866 VSS VDD  in_valid n713 n715 NAND2xp33_ASAP7_75t_R
XU867 VSS VDD  in_valid n194 n714 OR2x2_ASAP7_75t_R
XU868 VSS VDD  n537 n718 n589 n757 MAJIxp5_ASAP7_75t_R
XU869 VSS VDD  n212 n757 n719 XOR2xp5_ASAP7_75t_R
XU870 VSS VDD  n194 n719 A5  n720 HAxp5_ASAP7_75t_R
XU871 VSS VDD  in_valid n720 n722 NAND2xp33_ASAP7_75t_R
XU872 VSS VDD  Out_OFM[2] n395 n721 NAND2xp33_ASAP7_75t_R
XU873 VSS VDD  n723 n278 n262 n767 MAJIxp5_ASAP7_75t_R
XU874 VSS VDD  n767 n808 A6  n724 HAxp5_ASAP7_75t_R
XU875 VSS VDD  in_valid n725 n727 NAND2xp33_ASAP7_75t_R
XU876 VSS VDD  n774 n390 n726 NAND2xp33_ASAP7_75t_R
XU877 VSS VDD  n728 n246 n230 n762 MAJIxp5_ASAP7_75t_R
XU878 VSS VDD  n762 n830 A7  n729 HAxp5_ASAP7_75t_R
XU879 VSS VDD  in_valid n730 n732 NAND2xp33_ASAP7_75t_R
XU880 VSS VDD  n382 n574 n731 NAND2xp33_ASAP7_75t_R
XU881 VSS VDD  n544 n540 n805 NAND2xp33_ASAP7_75t_R
XU882 VSS VDD  n316 n348 n735 NOR2xp33_ASAP7_75t_R
XU883 VSS VDD  n346 n318 n733 NOR2xp33_ASAP7_75t_R
XU884 VSS VDD  n735 n733 A8  n804 HAxp5_ASAP7_75t_R
XU885 VSS VDD  n805 n804 n803 A9  n736 FAx1_ASAP7_75t_R
XU886 VSS VDD  in_valid n736 n738 NAND2xp33_ASAP7_75t_R
XU887 VSS VDD  in_valid n278 n737 OR2x2_ASAP7_75t_R
XU888 VSS VDD  n563 n547 n794 NAND2xp33_ASAP7_75t_R
XU889 VSS VDD  n292 n324 n741 NOR2xp33_ASAP7_75t_R
XU890 VSS VDD  n322 n294 n739 NOR2xp33_ASAP7_75t_R
XU891 VSS VDD  n741 n739 A10  n793 HAxp5_ASAP7_75t_R
XU892 VSS VDD  n794 n793 n792 A11  n742 FAx1_ASAP7_75t_R
XU893 VSS VDD  in_valid n742 n744 NAND2xp33_ASAP7_75t_R
XU894 VSS VDD  in_valid n230 n743 OR2x2_ASAP7_75t_R
XU895 VSS VDD  n564 n549 n827 NAND2xp33_ASAP7_75t_R
XU896 VSS VDD  n300 n332 n747 NOR2xp33_ASAP7_75t_R
XU897 VSS VDD  n330 n302 n745 NOR2xp33_ASAP7_75t_R
XU898 VSS VDD  n747 n745 A12  n826 HAxp5_ASAP7_75t_R
XU899 VSS VDD  n827 n826 n825 A13  n748 FAx1_ASAP7_75t_R
XU900 VSS VDD  in_valid n748 n750 NAND2xp33_ASAP7_75t_R
XU901 VSS VDD  in_valid n246 n749 OR2x2_ASAP7_75t_R
XU902 VSS VDD  n555 n538 n816 NAND2xp33_ASAP7_75t_R
XU903 VSS VDD  n308 n340 n753 NOR2xp33_ASAP7_75t_R
XU904 VSS VDD  n338 n310 n751 NOR2xp33_ASAP7_75t_R
XU905 VSS VDD  n753 n751 A14  n815 HAxp5_ASAP7_75t_R
XU906 VSS VDD  n816 n815 n814 A15  n754 FAx1_ASAP7_75t_R
XU907 VSS VDD  in_valid n754 n756 NAND2xp33_ASAP7_75t_R
XU908 VSS VDD  in_valid n262 n755 OR2x2_ASAP7_75t_R
XU909 VSS VDD  n212 n757 n194 n773 MAJIxp5_ASAP7_75t_R
XU910 VSS VDD  n773 n571 A16  n758 HAxp5_ASAP7_75t_R
XU911 VSS VDD  n758 n772 A17  n759 HAxp5_ASAP7_75t_R
XU912 VSS VDD  in_valid n759 n761 NAND2xp33_ASAP7_75t_R
XU913 VSS VDD  Out_OFM[3] n433 n760 NAND2xp33_ASAP7_75t_R
XU914 VSS VDD  n578 n762 n797 n779 MAJIxp5_ASAP7_75t_R
XU915 VSS VDD  n779 n250 n763 XOR2xp5_ASAP7_75t_R
XU916 VSS VDD  n234 n763 A18  n764 HAxp5_ASAP7_75t_R
XU917 VSS VDD  in_valid n764 n766 NAND2xp33_ASAP7_75t_R
XU918 VSS VDD  in_valid n198 n765 OR2x2_ASAP7_75t_R
XU919 VSS VDD  n576 n767 n819 n784 MAJIxp5_ASAP7_75t_R
XU920 VSS VDD  n784 n282 n768 XOR2xp5_ASAP7_75t_R
XU921 VSS VDD  n266 n768 A19  n769 HAxp5_ASAP7_75t_R
XU922 VSS VDD  in_valid n769 n771 NAND2xp33_ASAP7_75t_R
XU923 VSS VDD  in_valid n216 n770 OR2x2_ASAP7_75t_R
XU924 VSS VDD  n774 n773 n574 n871 MAJIxp5_ASAP7_75t_R
XU925 VSS VDD  n216 n871 n775 XOR2xp5_ASAP7_75t_R
XU926 VSS VDD  n198 n775 A20  n776 HAxp5_ASAP7_75t_R
XU927 VSS VDD  in_valid n776 n778 NAND2xp33_ASAP7_75t_R
XU928 VSS VDD  Out_OFM[4] n402 n777 NAND2xp33_ASAP7_75t_R
XU929 VSS VDD  n779 n250 n234 n833 MAJIxp5_ASAP7_75t_R
XU930 VSS VDD  n833 n904 A21  n780 HAxp5_ASAP7_75t_R
XU931 VSS VDD  in_valid n781 n783 NAND2xp33_ASAP7_75t_R
XU932 VSS VDD  n573 n403 n782 NAND2xp33_ASAP7_75t_R
XU933 VSS VDD  n784 n282 n266 n837 MAJIxp5_ASAP7_75t_R
XU934 VSS VDD  n837 n898 A22  n785 HAxp5_ASAP7_75t_R
XU935 VSS VDD  in_valid n786 n788 NAND2xp33_ASAP7_75t_R
XU936 VSS VDD  n890 n394 n787 NAND2xp33_ASAP7_75t_R
XU937 VSS VDD  n292 n548 n425 n588 mult_x_4_n36 NOR4xp25_ASAP7_75t_R
XU938 VSS VDD  n425 n292 n790 NOR2xp33_ASAP7_75t_R
XU939 VSS VDD  n548 n588 n789 NOR2xp33_ASAP7_75t_R
XU940 VSS VDD  n790 n789 n791 NOR2xp33_ASAP7_75t_R
XU941 VSS VDD  n794 n793 n792 n856 MAJIxp5_ASAP7_75t_R
XU942 VSS VDD  n856 n423 A23  n795 HAxp5_ASAP7_75t_R
XU943 VSS VDD  n857 n795 A24  n796 HAxp5_ASAP7_75t_R
XU944 VSS VDD  in_valid n796 n799 NAND2xp33_ASAP7_75t_R
XU945 VSS VDD  n797 n393 n798 NAND2xp33_ASAP7_75t_R
XU946 VSS VDD  n316 n541 n428 n585 mult_x_1_n36 NOR4xp25_ASAP7_75t_R
XU947 VSS VDD  n428 n316 n801 NOR2xp33_ASAP7_75t_R
XU948 VSS VDD  n541 n585 n800 NOR2xp33_ASAP7_75t_R
XU949 VSS VDD  n801 n800 n802 NOR2xp33_ASAP7_75t_R
XU950 VSS VDD  n805 n804 n803 n861 MAJIxp5_ASAP7_75t_R
XU951 VSS VDD  n861 n422 A25  n806 HAxp5_ASAP7_75t_R
XU952 VSS VDD  n862 n806 A26  n807 HAxp5_ASAP7_75t_R
XU953 VSS VDD  in_valid n807 n810 NAND2xp33_ASAP7_75t_R
XU954 VSS VDD  n576 n419 n809 NAND2xp33_ASAP7_75t_R
XU955 VSS VDD  n308 n539 n429 n586 mult_x_2_n36 NOR4xp25_ASAP7_75t_R
XU956 VSS VDD  n429 n308 n812 NOR2xp33_ASAP7_75t_R
XU957 VSS VDD  n539 n586 n811 NOR2xp33_ASAP7_75t_R
XU958 VSS VDD  n812 n811 n813 NOR2xp33_ASAP7_75t_R
XU959 VSS VDD  n816 n815 n814 n866 MAJIxp5_ASAP7_75t_R
XU960 VSS VDD  n866 n421 A27  n817 HAxp5_ASAP7_75t_R
XU961 VSS VDD  n867 n817 A28  n818 HAxp5_ASAP7_75t_R
XU962 VSS VDD  in_valid n818 n821 NAND2xp33_ASAP7_75t_R
XU963 VSS VDD  n819 n406 n820 NAND2xp33_ASAP7_75t_R
XU964 VSS VDD  n300 n550 n427 n587 mult_x_3_n36 NOR4xp25_ASAP7_75t_R
XU965 VSS VDD  n427 n300 n823 NOR2xp33_ASAP7_75t_R
XU966 VSS VDD  n550 n587 n822 NOR2xp33_ASAP7_75t_R
XU967 VSS VDD  n823 n822 n824 NOR2xp33_ASAP7_75t_R
XU968 VSS VDD  n827 n826 n825 n851 MAJIxp5_ASAP7_75t_R
XU969 VSS VDD  n851 n424 A29  n828 HAxp5_ASAP7_75t_R
XU970 VSS VDD  n852 n828 A30  n829 HAxp5_ASAP7_75t_R
XU971 VSS VDD  in_valid n829 n832 NAND2xp33_ASAP7_75t_R
XU972 VSS VDD  n578 n441 n831 NAND2xp33_ASAP7_75t_R
XU973 VSS VDD  n577 n833 n916 n846 MAJIxp5_ASAP7_75t_R
XU974 VSS VDD  n580 n240 n508 n834 MAJIxp5_ASAP7_75t_R
XU975 VSS VDD  in_valid n834 n836 NAND2xp33_ASAP7_75t_R
XU976 VSS VDD  n206 in_valid n835 OR2x2_ASAP7_75t_R
XU977 VSS VDD  n575 n837 n910 n841 MAJIxp5_ASAP7_75t_R
XU978 VSS VDD  n579 n272 n509 n838 MAJIxp5_ASAP7_75t_R
XU979 VSS VDD  in_valid n838 n840 NAND2xp33_ASAP7_75t_R
XU980 VSS VDD  n224 in_valid n839 OR2x2_ASAP7_75t_R
XU981 VSS VDD  n841 n286 n842 XOR2xp5_ASAP7_75t_R
XU982 VSS VDD  n270 n842 A31  n843 HAxp5_ASAP7_75t_R
XU983 VSS VDD  in_valid n843 n845 NAND2xp33_ASAP7_75t_R
XU984 VSS VDD  in_valid n220 n844 OR2x2_ASAP7_75t_R
XU985 VSS VDD  n846 n254 n847 XOR2xp5_ASAP7_75t_R
XU986 VSS VDD  n238 n847 A32  n848 HAxp5_ASAP7_75t_R
XU987 VSS VDD  in_valid n848 n850 NAND2xp33_ASAP7_75t_R
XU988 VSS VDD  in_valid n202 n849 OR2x2_ASAP7_75t_R
XU989 VSS VDD  n424 n852 n851 n901 MAJIxp5_ASAP7_75t_R
XU990 VSS VDD  mult_x_3_n30 n901 mult_x_3_n34 A33  n853 FAx1_ASAP7_75t_R
XU991 VSS VDD  in_valid n853 n855 NAND2xp33_ASAP7_75t_R
XU992 VSS VDD  n250 in_valid n854 OR2x2_ASAP7_75t_R
XU993 VSS VDD  n423 n857 n856 n913 MAJIxp5_ASAP7_75t_R
XU994 VSS VDD  mult_x_4_n30 n913 mult_x_4_n34 A34  n858 FAx1_ASAP7_75t_R
XU995 VSS VDD  in_valid n858 n860 NAND2xp33_ASAP7_75t_R
XU996 VSS VDD  n234 in_valid n859 OR2x2_ASAP7_75t_R
XU997 VSS VDD  n422 n862 n861 n895 MAJIxp5_ASAP7_75t_R
XU998 VSS VDD  mult_x_1_n30 n895 mult_x_1_n34 A35  n863 FAx1_ASAP7_75t_R
XU999 VSS VDD  in_valid n863 n865 NAND2xp33_ASAP7_75t_R
XU1000 VSS VDD  n282 in_valid n864 OR2x2_ASAP7_75t_R
XU1001 VSS VDD  n421 n867 n866 n907 MAJIxp5_ASAP7_75t_R
XU1002 VSS VDD  mult_x_2_n30 n907 mult_x_2_n34 A36  n868 FAx1_ASAP7_75t_R
XU1003 VSS VDD  in_valid n868 n870 NAND2xp33_ASAP7_75t_R
XU1004 VSS VDD  n266 in_valid n869 OR2x2_ASAP7_75t_R
XU1005 VSS VDD  n216 n871 n198 n889 MAJIxp5_ASAP7_75t_R
XU1006 VSS VDD  n889 n570 A37  n872 HAxp5_ASAP7_75t_R
XU1007 VSS VDD  n872 n888 A38  n873 HAxp5_ASAP7_75t_R
XU1008 VSS VDD  in_valid n873 n875 NAND2xp33_ASAP7_75t_R
XU1009 VSS VDD  Out_OFM[5] n407 n874 NAND2xp33_ASAP7_75t_R
XU1010 VSS VDD  n921 n388 n881 NAND2xp33_ASAP7_75t_R
XU1011 VSS VDD  n944 n447 n877 NAND2xp33_ASAP7_75t_R
XU1012 VSS VDD  n579 n509 n876 NAND2xp33_ASAP7_75t_R
XU1013 VSS VDD  n878 n272 n879 XOR2xp5_ASAP7_75t_R
XU1014 VSS VDD  in_valid n879 n880 NAND2xp33_ASAP7_75t_R
XU1015 VSS VDD  n572 n415 n887 NAND2xp33_ASAP7_75t_R
XU1016 VSS VDD  n938 n446 n883 NAND2xp33_ASAP7_75t_R
XU1017 VSS VDD  n580 n508 n882 NAND2xp33_ASAP7_75t_R
XU1018 VSS VDD  n884 n240 n885 XOR2xp5_ASAP7_75t_R
XU1019 VSS VDD  in_valid n885 n886 NAND2xp33_ASAP7_75t_R
XU1020 VSS VDD  n890 n889 n573 n919 MAJIxp5_ASAP7_75t_R
XU1021 VSS VDD  n220 n919 n891 XOR2xp5_ASAP7_75t_R
XU1022 VSS VDD  n202 n891 A39  n892 HAxp5_ASAP7_75t_R
XU1023 VSS VDD  in_valid n892 n894 NAND2xp33_ASAP7_75t_R
XU1024 VSS VDD  Out_OFM[6] n401 n893 NAND2xp33_ASAP7_75t_R
XU1025 VSS VDD  mult_x_1_n29 n442 A40  n896 HAxp5_ASAP7_75t_R
XU1026 VSS VDD  mult_x_1_n26 n896 A41  n897 HAxp5_ASAP7_75t_R
XU1027 VSS VDD  in_valid n897 n900 NAND2xp33_ASAP7_75t_R
XU1028 VSS VDD  n575 n435 n899 NAND2xp33_ASAP7_75t_R
XU1029 VSS VDD  mult_x_3_n29 n443 A42  n902 HAxp5_ASAP7_75t_R
XU1030 VSS VDD  mult_x_3_n26 n902 A43  n903 HAxp5_ASAP7_75t_R
XU1031 VSS VDD  in_valid n903 n906 NAND2xp33_ASAP7_75t_R
XU1032 VSS VDD  n577 n408 n905 NAND2xp33_ASAP7_75t_R
XU1033 VSS VDD  mult_x_2_n29 n444 A44  n908 HAxp5_ASAP7_75t_R
XU1034 VSS VDD  mult_x_2_n26 n908 A45  n909 HAxp5_ASAP7_75t_R
XU1035 VSS VDD  in_valid n909 n912 NAND2xp33_ASAP7_75t_R
XU1036 VSS VDD  n910 n391 n911 NAND2xp33_ASAP7_75t_R
XU1037 VSS VDD  mult_x_4_n29 n445 A46  n914 HAxp5_ASAP7_75t_R
XU1038 VSS VDD  mult_x_4_n26 n914 A47  n915 HAxp5_ASAP7_75t_R
XU1039 VSS VDD  in_valid n915 n918 NAND2xp33_ASAP7_75t_R
XU1040 VSS VDD  n916 n420 n917 NAND2xp33_ASAP7_75t_R
XU1041 VSS VDD  n220 n919 n202 n947 MAJIxp5_ASAP7_75t_R
XU1042 VSS VDD  n921 n947 n572 n972 MAJIxp5_ASAP7_75t_R
XU1043 VSS VDD  n206 n224 n972 n922 MAJIxp5_ASAP7_75t_R
XU1044 VSS VDD  in_valid n922 n924 NAND2xp33_ASAP7_75t_R
XU1045 VSS VDD  Out_OFM[9] n432 n923 NAND2xp33_ASAP7_75t_R
XU1046 VSS VDD  n925 mult_x_4_n29 mult_x_4_n26 n958 MAJx2_ASAP7_75t_R
XU1047 VSS VDD  n560 n926 n957 NAND2xp33_ASAP7_75t_R
XU1048 VSS VDD  mult_x_4_n25 n958 n957 n927 MAJIxp5_ASAP7_75t_R
XU1049 VSS VDD  in_valid n927 n929 NAND2xp33_ASAP7_75t_R
XU1050 VSS VDD  n240 in_valid n928 OR2x2_ASAP7_75t_R
XU1051 VSS VDD  n930 mult_x_2_n29 mult_x_2_n26 n968 MAJx2_ASAP7_75t_R
XU1052 VSS VDD  n545 n931 n967 NAND2xp33_ASAP7_75t_R
XU1053 VSS VDD  mult_x_2_n25 n968 n967 n932 MAJIxp5_ASAP7_75t_R
XU1054 VSS VDD  in_valid n932 n934 NAND2xp33_ASAP7_75t_R
XU1055 VSS VDD  n272 in_valid n933 OR2x2_ASAP7_75t_R
XU1056 VSS VDD  n935 mult_x_3_n29 mult_x_3_n26 n953 MAJx2_ASAP7_75t_R
XU1057 VSS VDD  n561 n936 n952 NAND2xp33_ASAP7_75t_R
XU1058 VSS VDD  mult_x_3_n25 n953 n952 n937 MAJIxp5_ASAP7_75t_R
XU1059 VSS VDD  in_valid n937 n940 NAND2xp33_ASAP7_75t_R
XU1060 VSS VDD  n938 n414 n939 NAND2xp33_ASAP7_75t_R
XU1061 VSS VDD  n941 mult_x_1_n29 mult_x_1_n26 n963 MAJx2_ASAP7_75t_R
XU1062 VSS VDD  n562 n942 n962 NAND2xp33_ASAP7_75t_R
XU1063 VSS VDD  mult_x_1_n25 n963 n962 n943 MAJIxp5_ASAP7_75t_R
XU1064 VSS VDD  in_valid n943 n946 NAND2xp33_ASAP7_75t_R
XU1065 VSS VDD  n944 n392 n945 NAND2xp33_ASAP7_75t_R
XU1066 VSS VDD  n947 n569 A48  n948 HAxp5_ASAP7_75t_R
XU1067 VSS VDD  n948 n920 A49  n949 HAxp5_ASAP7_75t_R
XU1068 VSS VDD  in_valid n949 n951 NAND2xp33_ASAP7_75t_R
XU1069 VSS VDD  Out_OFM[7] n410 n950 NAND2xp33_ASAP7_75t_R
XU1070 VSS VDD  mult_x_3_n25 n953 n952 A50  n954 FAx1_ASAP7_75t_R
XU1071 VSS VDD  in_valid n954 n956 NAND2xp33_ASAP7_75t_R
XU1072 VSS VDD  n254 in_valid n955 OR2x2_ASAP7_75t_R
XU1073 VSS VDD  mult_x_4_n25 n958 n957 A51  n959 FAx1_ASAP7_75t_R
XU1074 VSS VDD  in_valid n959 n961 NAND2xp33_ASAP7_75t_R
XU1075 VSS VDD  n238 in_valid n960 OR2x2_ASAP7_75t_R
XU1076 VSS VDD  mult_x_1_n25 n963 n962 A52  n964 FAx1_ASAP7_75t_R
XU1077 VSS VDD  in_valid n964 n966 NAND2xp33_ASAP7_75t_R
XU1078 VSS VDD  n286 in_valid n965 OR2x2_ASAP7_75t_R
XU1079 VSS VDD  mult_x_2_n25 n968 n967 A53  n969 FAx1_ASAP7_75t_R
XU1080 VSS VDD  in_valid n969 n971 NAND2xp33_ASAP7_75t_R
XU1081 VSS VDD  n270 in_valid n970 OR2x2_ASAP7_75t_R
XU1082 VSS VDD  n224 n972 n974 NOR2xp33_ASAP7_75t_R
XU1083 VSS VDD  n224 n972 n973 AND2x2_ASAP7_75t_R
XU1084 VSS VDD  n206 n975 A54  n976 HAxp5_ASAP7_75t_R
XU1085 VSS VDD  in_valid n976 n978 NAND2xp33_ASAP7_75t_R
XU1086 VSS VDD  Out_OFM[8] n440 n977 NAND2xp33_ASAP7_75t_R
XU1087 VSS VDD  n316 n431 n585 n348 mult_x_1_n31 NOR4xp25_ASAP7_75t_R
XU1088 VSS VDD  n431 n348 n980 NOR2xp33_ASAP7_75t_R
XU1089 VSS VDD  n585 n316 n979 NOR2xp33_ASAP7_75t_R
XU1090 VSS VDD  n980 n979 n981 NOR2xp33_ASAP7_75t_R
XU1091 VSS VDD  mult_x_1_n31 n981 mult_x_1_n32 NOR2xp33_ASAP7_75t_R
XU1092 VSS VDD  n316 n348 n346 n318 mult_x_1_n38 NOR4xp25_ASAP7_75t_R
XU1093 VSS VDD  n585 n318 mult_x_1_n41 NOR2xp33_ASAP7_75t_R
XU1094 VSS VDD  n431 n428 mult_x_1_n44 NOR2xp33_ASAP7_75t_R
XU1095 VSS VDD  n428 n318 mult_x_1_n45 NOR2xp33_ASAP7_75t_R
XU1096 VSS VDD  n348 n318 mult_x_1_n49 NOR2xp33_ASAP7_75t_R
XU1097 VSS VDD  n431 n346 mult_x_1_n52 NOR2xp33_ASAP7_75t_R
XU1098 VSS VDD  n308 n546 n586 n340 mult_x_2_n31 NOR4xp25_ASAP7_75t_R
XU1099 VSS VDD  n546 n340 n983 NOR2xp33_ASAP7_75t_R
XU1100 VSS VDD  n586 n308 n982 NOR2xp33_ASAP7_75t_R
XU1101 VSS VDD  n983 n982 n984 NOR2xp33_ASAP7_75t_R
XU1102 VSS VDD  mult_x_2_n31 n984 mult_x_2_n32 NOR2xp33_ASAP7_75t_R
XU1103 VSS VDD  n308 n340 n338 n310 mult_x_2_n38 NOR4xp25_ASAP7_75t_R
XU1104 VSS VDD  n586 n310 mult_x_2_n41 NOR2xp33_ASAP7_75t_R
XU1105 VSS VDD  n546 n429 mult_x_2_n44 NOR2xp33_ASAP7_75t_R
XU1106 VSS VDD  n429 n310 mult_x_2_n45 NOR2xp33_ASAP7_75t_R
XU1107 VSS VDD  n340 n310 mult_x_2_n49 NOR2xp33_ASAP7_75t_R
XU1108 VSS VDD  n546 n338 mult_x_2_n52 NOR2xp33_ASAP7_75t_R
XU1109 VSS VDD  n300 n426 n587 n332 mult_x_3_n31 NOR4xp25_ASAP7_75t_R
XU1110 VSS VDD  n426 n332 n986 NOR2xp33_ASAP7_75t_R
XU1111 VSS VDD  n587 n300 n985 NOR2xp33_ASAP7_75t_R
XU1112 VSS VDD  n986 n985 n987 NOR2xp33_ASAP7_75t_R
XU1113 VSS VDD  mult_x_3_n31 n987 mult_x_3_n32 NOR2xp33_ASAP7_75t_R
XU1114 VSS VDD  n300 n332 n330 n302 mult_x_3_n38 NOR4xp25_ASAP7_75t_R
XU1115 VSS VDD  n587 n302 mult_x_3_n41 NOR2xp33_ASAP7_75t_R
XU1116 VSS VDD  n426 n427 mult_x_3_n44 NOR2xp33_ASAP7_75t_R
XU1117 VSS VDD  n427 n302 mult_x_3_n45 NOR2xp33_ASAP7_75t_R
XU1118 VSS VDD  n332 n302 mult_x_3_n49 NOR2xp33_ASAP7_75t_R
XU1119 VSS VDD  n426 n330 mult_x_3_n52 NOR2xp33_ASAP7_75t_R
XU1120 VSS VDD  n292 n430 n588 n324 mult_x_4_n31 NOR4xp25_ASAP7_75t_R
XU1121 VSS VDD  n430 n324 n989 NOR2xp33_ASAP7_75t_R
XU1122 VSS VDD  n588 n292 n988 NOR2xp33_ASAP7_75t_R
XU1123 VSS VDD  n989 n988 n990 NOR2xp33_ASAP7_75t_R
XU1124 VSS VDD  mult_x_4_n31 n990 mult_x_4_n32 NOR2xp33_ASAP7_75t_R
XU1125 VSS VDD  n292 n324 n322 n294 mult_x_4_n38 NOR4xp25_ASAP7_75t_R
XU1126 VSS VDD  n588 n294 mult_x_4_n41 NOR2xp33_ASAP7_75t_R
XU1127 VSS VDD  n430 n425 mult_x_4_n44 NOR2xp33_ASAP7_75t_R
XU1128 VSS VDD  n425 n294 mult_x_4_n45 NOR2xp33_ASAP7_75t_R
XU1129 VSS VDD  n324 n294 mult_x_4_n49 NOR2xp33_ASAP7_75t_R
XU1130 VSS VDD  n430 n322 mult_x_4_n52 NOR2xp33_ASAP7_75t_R
.ENDS


